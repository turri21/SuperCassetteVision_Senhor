    ird_lut['h00a] = {UA_MOV_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h00b] = {UA_MOV_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h00c] = {UA_MOV_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h00d] = {UA_MOV_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h00e] = {UA_MOV_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h00f] = {UA_MOV_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h01a] = {UA_MOV_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h01b] = {UA_MOV_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h01c] = {UA_MOV_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h01d] = {UA_MOV_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h01e] = {UA_MOV_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h01f] = {UA_MOV_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h068] = {UA_MOV_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h069] = {UA_MOV_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h06a] = {UA_MOV_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h06b] = {UA_MOV_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h06c] = {UA_MOV_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h06d] = {UA_MOV_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h06e] = {UA_MOV_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h069] = {UA_MOV_RF_IR210_IMM_L1, 1'd0, 2'd1, ISEFM_L1};
    ird_lut['h06f] = {UA_MOV_RF_IR210_IMM_L0, 1'd0, 2'd1, ISEFM_L0};
    ird_lut['h028] = {UA_LD_A_WA, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h004] = {UA_LDX_SP_IMM, 1'd0, 2'd2, ISEFM_NONE};
    ird_lut['h014] = {UA_LDX_BC_IMM, 1'd0, 2'd2, ISEFM_NONE};
    ird_lut['h024] = {UA_LDX_DE_IMM, 1'd0, 2'd2, ISEFM_NONE};
    ird_lut['h034] = {UA_LDX_HL_IMM_L0, 1'd0, 2'd2, ISEFM_L0};
    ird_lut['h029] = {UA_LDAX, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h02a] = {UA_LDAX, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h02b] = {UA_LDAX, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h02c] = {UA_LDAX, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h02d] = {UA_LDAX, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h02e] = {UA_LDAX, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h02f] = {UA_LDAX, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h039] = {UA_STX_A, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h03a] = {UA_STX_A, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h03b] = {UA_STX_A, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h03c] = {UA_STX_A, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h03d] = {UA_STX_A, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h03e] = {UA_STX_A, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h03f] = {UA_STX_A, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h049] = {UA_STX_RF_W, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h04a] = {UA_STX_RF_W, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h04b] = {UA_STX_RF_W, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h038] = {UA_STW_A, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h071] = {UA_STW_IMM, 1'd0, 2'd2, ISEFM_NONE};
    ird_lut['h021] = {UA_TABLE, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h031] = {UA_BLOCK, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h010] = {UA_EX, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h011] = {UA_EXX, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h005] = {UA_AND_WA_IMM, 1'd0, 2'd2, ISEFM_NONE};
    ird_lut['h015] = {UA_OR_WA_IMM, 1'd0, 2'd2, ISEFM_NONE};
    ird_lut['h007] = {UA_AND_A_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h016] = {UA_XOR_A_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h017] = {UA_OR_A_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h025] = {UA_CMPBNB_WA_IMM, 1'd0, 2'd2, ISEFM_NONE};
    ird_lut['h035] = {UA_CMPB_WA_IMM, 1'd0, 2'd2, ISEFM_NONE};
    ird_lut['h045] = {UA_BITNZ_WA_IMM, 1'd0, 2'd2, ISEFM_NONE};
    ird_lut['h055] = {UA_BITZ_WA_IMM, 1'd0, 2'd2, ISEFM_NONE};
    ird_lut['h065] = {UA_CMPNZ_WA_IMM, 1'd0, 2'd2, ISEFM_NONE};
    ird_lut['h075] = {UA_CMPZ_WA_IMM, 1'd0, 2'd2, ISEFM_NONE};
    ird_lut['h027] = {UA_CMPBNB_A_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h037] = {UA_CMPB_A_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h047] = {UA_BITNZ_A_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h057] = {UA_BITZ_A_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h067] = {UA_CMPNZ_A_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h077] = {UA_CMPZ_A_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h026] = {UA_ADDNC_A_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h036] = {UA_SUBNB_A_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h046] = {UA_ADD_A_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h056] = {UA_ADC_A_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h066] = {UA_SUB_A_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h076] = {UA_SBB_A_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h020] = {UA_INCR_WA, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h030] = {UA_DECR_WA, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h041] = {UA_INCR_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h042] = {UA_INCR_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h043] = {UA_INCR_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h051] = {UA_DECR_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h052] = {UA_DECR_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h053] = {UA_DECR_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h002] = {UA_INC_SP, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h012] = {UA_INC_BC, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h022] = {UA_INC_DE, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h032] = {UA_INC_HL, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h003] = {UA_DEC_SP, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h013] = {UA_DEC_BC, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h023] = {UA_DEC_DE, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h033] = {UA_DEC_HL, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h061] = {UA_DAA, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h0c0] = {UA_JR, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0c1] = {UA_JR, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0c2] = {UA_JR, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0c3] = {UA_JR, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0c4] = {UA_JR, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0c5] = {UA_JR, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0c6] = {UA_JR, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0c7] = {UA_JR, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0c8] = {UA_JR, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0c9] = {UA_JR, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0ca] = {UA_JR, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0cb] = {UA_JR, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0cc] = {UA_JR, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0cd] = {UA_JR, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0ce] = {UA_JR, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0cf] = {UA_JR, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0d0] = {UA_JR, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0d1] = {UA_JR, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0d2] = {UA_JR, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0d3] = {UA_JR, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0d4] = {UA_JR, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0d5] = {UA_JR, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0d6] = {UA_JR, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0d7] = {UA_JR, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0d8] = {UA_JR, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0d9] = {UA_JR, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0da] = {UA_JR, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0db] = {UA_JR, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0dc] = {UA_JR, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0dd] = {UA_JR, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0de] = {UA_JR, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0df] = {UA_JR, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0e0] = {UA_JR, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0e1] = {UA_JR, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0e2] = {UA_JR, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0e3] = {UA_JR, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0e4] = {UA_JR, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0e5] = {UA_JR, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0e6] = {UA_JR, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0e7] = {UA_JR, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0e8] = {UA_JR, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0e9] = {UA_JR, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0ea] = {UA_JR, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0eb] = {UA_JR, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0ec] = {UA_JR, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0ed] = {UA_JR, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0ee] = {UA_JR, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0ef] = {UA_JR, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0f0] = {UA_JR, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0f1] = {UA_JR, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0f2] = {UA_JR, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0f3] = {UA_JR, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0f4] = {UA_JR, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0f5] = {UA_JR, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0f6] = {UA_JR, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0f7] = {UA_JR, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0f8] = {UA_JR, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0f9] = {UA_JR, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0fa] = {UA_JR, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0fb] = {UA_JR, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0fc] = {UA_JR, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0fd] = {UA_JR, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0fe] = {UA_JR, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0ff] = {UA_JR, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h04e] = {UA_JRE_P, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h04f] = {UA_JRE_N, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h054] = {UA_JMP, 1'd0, 2'd2, ISEFM_NONE};
    ird_lut['h073] = {UA_JB, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h044] = {UA_CALL, 1'd0, 2'd2, ISEFM_NONE};
    ird_lut['h063] = {UA_CALB, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h078] = {UA_CALF, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h079] = {UA_CALF, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h07a] = {UA_CALF, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h07b] = {UA_CALF, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h07c] = {UA_CALF, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h07d] = {UA_CALF, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h07e] = {UA_CALF, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h07f] = {UA_CALF, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h080] = {UA_CALT, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h081] = {UA_CALT, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h082] = {UA_CALT, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h083] = {UA_CALT, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h084] = {UA_CALT, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h085] = {UA_CALT, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h086] = {UA_CALT, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h087] = {UA_CALT, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h088] = {UA_CALT, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h089] = {UA_CALT, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h08a] = {UA_CALT, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h08b] = {UA_CALT, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h08c] = {UA_CALT, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h08d] = {UA_CALT, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h08e] = {UA_CALT, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h08f] = {UA_CALT, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h090] = {UA_CALT, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h091] = {UA_CALT, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h092] = {UA_CALT, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h093] = {UA_CALT, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h094] = {UA_CALT, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h095] = {UA_CALT, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h096] = {UA_CALT, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h097] = {UA_CALT, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h098] = {UA_CALT, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h099] = {UA_CALT, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h09a] = {UA_CALT, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h09b] = {UA_CALT, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h09c] = {UA_CALT, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h09d] = {UA_CALT, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h09e] = {UA_CALT, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h09f] = {UA_CALT, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0a0] = {UA_CALT, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0a1] = {UA_CALT, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0a2] = {UA_CALT, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0a3] = {UA_CALT, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0a4] = {UA_CALT, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0a5] = {UA_CALT, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0a6] = {UA_CALT, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0a7] = {UA_CALT, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0a8] = {UA_CALT, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0a9] = {UA_CALT, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0aa] = {UA_CALT, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0ab] = {UA_CALT, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0ac] = {UA_CALT, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0ad] = {UA_CALT, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0ae] = {UA_CALT, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0af] = {UA_CALT, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0b0] = {UA_CALT, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0b1] = {UA_CALT, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0b2] = {UA_CALT, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0b3] = {UA_CALT, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0b4] = {UA_CALT, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0b5] = {UA_CALT, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0b6] = {UA_CALT, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0b7] = {UA_CALT, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0b8] = {UA_CALT, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0b9] = {UA_CALT, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0ba] = {UA_CALT, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0bb] = {UA_CALT, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0bc] = {UA_CALT, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0bd] = {UA_CALT, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0be] = {UA_CALT, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h0bf] = {UA_CALT, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h072] = {UA_INT, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h008] = {UA_RET, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h018] = {UA_RETS, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h062] = {UA_RETI, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h058] = {UA_BIT, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h059] = {UA_BIT, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h05a] = {UA_BIT, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h05b] = {UA_BIT, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h05c] = {UA_BIT, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h05d] = {UA_BIT, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h05e] = {UA_BIT, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h05f] = {UA_BIT, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h000] = {UA_NOP, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h019] = {UA_STM, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h130] = {UA_RLL_A_, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h131] = {UA_RLR_A_, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h132] = {UA_RLL_C_, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h133] = {UA_RLR_C_, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h134] = {UA_SLL_A_, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h135] = {UA_SLR_A_, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h136] = {UA_SLL_C_, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h137] = {UA_SLR_C_, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h10e] = {UA_PUSH_VA, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h10f] = {UA_POP_VA, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h11e] = {UA_PUSH_BC, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h11f] = {UA_POP_BC, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h12e] = {UA_PUSH_DE, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h12f] = {UA_POP_DE, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h13e] = {UA_PUSH_HL, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h13f] = {UA_POP_HL, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h100] = {UA_SKIP_I, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h101] = {UA_SKIP_I, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h102] = {UA_SKIP_I, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h103] = {UA_SKIP_I, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h104] = {UA_SKIP_I, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h10a] = {UA_SKIP_PSW_C, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h10c] = {UA_SKIP_PSW_Z, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h110] = {UA_SKIP_NI, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h111] = {UA_SKIP_NI, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h112] = {UA_SKIP_NI, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h113] = {UA_SKIP_NI, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h114] = {UA_SKIP_NI, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h11a] = {UA_SKIP_PSW_NC, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h11c] = {UA_SKIP_PSW_NZ, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h120] = {UA_EI, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h124] = {UA_DI, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h12a] = {UA_CLC, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h12b] = {UA_STC, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h138] = {UA_RLD, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h139] = {UA_RRD, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h2c0] = {UA_MOV_A_SPR_IR3, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h2c1] = {UA_MOV_A_SPR_IR3, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h2c2] = {UA_MOV_A_SPR_IR3, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h2c3] = {UA_MOV_A_SPR_IR3, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h2c4] = {UA_MOV_A_SPR_IR3, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h2c5] = {UA_MOV_A_SPR_IR3, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h2c6] = {UA_MOV_A_SPR_IR3, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h2c7] = {UA_MOV_A_SPR_IR3, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h2c8] = {UA_MOV_A_SPR_IR3, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h2c9] = {UA_MOV_A_SPR_IR3, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h3c0] = {UA_MOV_SPR_IR3_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h3c1] = {UA_MOV_SPR_IR3_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h3c2] = {UA_MOV_SPR_IR3_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h3c3] = {UA_MOV_SPR_IR3_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h3c4] = {UA_MOV_SPR_IR3_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h3c5] = {UA_MOV_SPR_IR3_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h3c6] = {UA_MOV_SPR_IR3_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h3c7] = {UA_MOV_SPR_IR3_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h3c8] = {UA_MOV_SPR_IR3_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h3c9] = {UA_MOV_SPR_IR3_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h420] = {UA_ADDNC_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h421] = {UA_ADDNC_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h422] = {UA_ADDNC_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h423] = {UA_ADDNC_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h424] = {UA_ADDNC_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h425] = {UA_ADDNC_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h426] = {UA_ADDNC_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h427] = {UA_ADDNC_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h430] = {UA_SUBNB_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h431] = {UA_SUBNB_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h432] = {UA_SUBNB_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h433] = {UA_SUBNB_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h434] = {UA_SUBNB_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h435] = {UA_SUBNB_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h436] = {UA_SUBNB_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h437] = {UA_SUBNB_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h440] = {UA_ADD_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h441] = {UA_ADD_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h442] = {UA_ADD_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h443] = {UA_ADD_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h444] = {UA_ADD_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h445] = {UA_ADD_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h446] = {UA_ADD_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h447] = {UA_ADD_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h450] = {UA_ADC_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h451] = {UA_ADC_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h452] = {UA_ADC_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h453] = {UA_ADC_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h454] = {UA_ADC_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h455] = {UA_ADC_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h456] = {UA_ADC_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h457] = {UA_ADC_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h460] = {UA_SUB_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h461] = {UA_SUB_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h462] = {UA_SUB_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h463] = {UA_SUB_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h464] = {UA_SUB_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h465] = {UA_SUB_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h466] = {UA_SUB_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h467] = {UA_SUB_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h470] = {UA_SBB_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h471] = {UA_SBB_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h472] = {UA_SBB_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h473] = {UA_SBB_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h474] = {UA_SBB_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h475] = {UA_SBB_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h476] = {UA_SBB_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h477] = {UA_SBB_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4a0] = {UA_ADDNC_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4a1] = {UA_ADDNC_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4a2] = {UA_ADDNC_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4a3] = {UA_ADDNC_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4a4] = {UA_ADDNC_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4a5] = {UA_ADDNC_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4a6] = {UA_ADDNC_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4a7] = {UA_ADDNC_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4b0] = {UA_SUBNB_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4b1] = {UA_SUBNB_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4b2] = {UA_SUBNB_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4b3] = {UA_SUBNB_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4b4] = {UA_SUBNB_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4b5] = {UA_SUBNB_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4b6] = {UA_SUBNB_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4b7] = {UA_SUBNB_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4c0] = {UA_ADD_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4c1] = {UA_ADD_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4c2] = {UA_ADD_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4c3] = {UA_ADD_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4c4] = {UA_ADD_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4c5] = {UA_ADD_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4c6] = {UA_ADD_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4c7] = {UA_ADD_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4d0] = {UA_ADC_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4d1] = {UA_ADC_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4d2] = {UA_ADC_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4d3] = {UA_ADC_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4d4] = {UA_ADC_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4d5] = {UA_ADC_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4d6] = {UA_ADC_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4d7] = {UA_ADC_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4e0] = {UA_SUB_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4e1] = {UA_SUB_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4e2] = {UA_SUB_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4e3] = {UA_SUB_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4e4] = {UA_SUB_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4e5] = {UA_SUB_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4e6] = {UA_SUB_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4e7] = {UA_SUB_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4f0] = {UA_SBB_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4f1] = {UA_SBB_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4f2] = {UA_SBB_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4f3] = {UA_SBB_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4f4] = {UA_SBB_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4f5] = {UA_SBB_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4f6] = {UA_SBB_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4f7] = {UA_SBB_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h408] = {UA_AND_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h409] = {UA_AND_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h40a] = {UA_AND_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h40b] = {UA_AND_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h40c] = {UA_AND_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h40d] = {UA_AND_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h40e] = {UA_AND_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h40f] = {UA_AND_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h410] = {UA_XOR_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h411] = {UA_XOR_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h412] = {UA_XOR_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h413] = {UA_XOR_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h414] = {UA_XOR_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h415] = {UA_XOR_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h416] = {UA_XOR_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h417] = {UA_XOR_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h418] = {UA_OR_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h419] = {UA_OR_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h41a] = {UA_OR_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h41b] = {UA_OR_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h41c] = {UA_OR_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h41d] = {UA_OR_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h41e] = {UA_OR_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h41f] = {UA_OR_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h488] = {UA_AND_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h489] = {UA_AND_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h48a] = {UA_AND_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h48b] = {UA_AND_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h48c] = {UA_AND_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h48d] = {UA_AND_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h48e] = {UA_AND_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h48f] = {UA_AND_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h490] = {UA_XOR_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h491] = {UA_XOR_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h492] = {UA_XOR_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h493] = {UA_XOR_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h494] = {UA_XOR_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h495] = {UA_XOR_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h496] = {UA_XOR_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h497] = {UA_XOR_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h498] = {UA_OR_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h499] = {UA_OR_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h49a] = {UA_OR_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h49b] = {UA_OR_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h49c] = {UA_OR_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h49d] = {UA_OR_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h49e] = {UA_OR_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h49f] = {UA_OR_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h428] = {UA_CMPBNB_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h429] = {UA_CMPBNB_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h42a] = {UA_CMPBNB_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h42b] = {UA_CMPBNB_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h42c] = {UA_CMPBNB_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h42d] = {UA_CMPBNB_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h42e] = {UA_CMPBNB_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h42f] = {UA_CMPBNB_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h438] = {UA_CMPB_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h439] = {UA_CMPB_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h43a] = {UA_CMPB_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h43b] = {UA_CMPB_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h43c] = {UA_CMPB_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h43d] = {UA_CMPB_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h43e] = {UA_CMPB_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h43f] = {UA_CMPB_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h468] = {UA_CMPNZ_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h469] = {UA_CMPNZ_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h46a] = {UA_CMPNZ_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h46b] = {UA_CMPNZ_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h46c] = {UA_CMPNZ_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h46d] = {UA_CMPNZ_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h46e] = {UA_CMPNZ_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h46f] = {UA_CMPNZ_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h478] = {UA_CMPZ_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h479] = {UA_CMPZ_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h47a] = {UA_CMPZ_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h47b] = {UA_CMPZ_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h47c] = {UA_CMPZ_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h47d] = {UA_CMPZ_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h47e] = {UA_CMPZ_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h47f] = {UA_CMPZ_RF_IR210_A, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4a8] = {UA_CMPBNB_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4a9] = {UA_CMPBNB_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4aa] = {UA_CMPBNB_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4ab] = {UA_CMPBNB_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4ac] = {UA_CMPBNB_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4ad] = {UA_CMPBNB_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4ae] = {UA_CMPBNB_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4af] = {UA_CMPBNB_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4b8] = {UA_CMPB_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4b9] = {UA_CMPB_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4ba] = {UA_CMPB_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4bb] = {UA_CMPB_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4bc] = {UA_CMPB_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4bd] = {UA_CMPB_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4be] = {UA_CMPB_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4bf] = {UA_CMPB_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4c8] = {UA_BITNZ_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4c9] = {UA_BITNZ_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4ca] = {UA_BITNZ_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4cb] = {UA_BITNZ_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4cc] = {UA_BITNZ_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4cd] = {UA_BITNZ_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4ce] = {UA_BITNZ_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4cf] = {UA_BITNZ_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4d8] = {UA_BITZ_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4d9] = {UA_BITZ_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4da] = {UA_BITZ_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4db] = {UA_BITZ_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4dc] = {UA_BITZ_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4dd] = {UA_BITZ_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4de] = {UA_BITZ_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4df] = {UA_BITZ_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4e8] = {UA_CMPNZ_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4e9] = {UA_CMPNZ_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4ea] = {UA_CMPNZ_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4eb] = {UA_CMPNZ_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4ec] = {UA_CMPNZ_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4ed] = {UA_CMPNZ_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4ee] = {UA_CMPNZ_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4ef] = {UA_CMPNZ_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4f8] = {UA_CMPZ_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4f9] = {UA_CMPZ_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4fa] = {UA_CMPZ_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4fb] = {UA_CMPZ_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4fc] = {UA_CMPZ_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4fd] = {UA_CMPZ_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4fe] = {UA_CMPZ_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h4ff] = {UA_CMPZ_A_RF_IR210, 1'd1, 2'd0, ISEFM_NONE};
    ird_lut['h520] = {UA_ADDNC_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h521] = {UA_ADDNC_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h522] = {UA_ADDNC_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h523] = {UA_ADDNC_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h524] = {UA_ADDNC_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h525] = {UA_ADDNC_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h526] = {UA_ADDNC_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h527] = {UA_ADDNC_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h530] = {UA_SUBNB_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h531] = {UA_SUBNB_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h532] = {UA_SUBNB_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h533] = {UA_SUBNB_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h534] = {UA_SUBNB_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h535] = {UA_SUBNB_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h536] = {UA_SUBNB_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h537] = {UA_SUBNB_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h540] = {UA_ADD_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h541] = {UA_ADD_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h542] = {UA_ADD_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h543] = {UA_ADD_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h544] = {UA_ADD_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h545] = {UA_ADD_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h546] = {UA_ADD_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h547] = {UA_ADD_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h550] = {UA_ADC_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h551] = {UA_ADC_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h552] = {UA_ADC_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h553] = {UA_ADC_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h554] = {UA_ADC_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h555] = {UA_ADC_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h556] = {UA_ADC_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h557] = {UA_ADC_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h560] = {UA_SUB_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h561] = {UA_SUB_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h562] = {UA_SUB_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h563] = {UA_SUB_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h564] = {UA_SUB_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h565] = {UA_SUB_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h566] = {UA_SUB_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h567] = {UA_SUB_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h570] = {UA_SBB_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h571] = {UA_SBB_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h572] = {UA_SBB_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h573] = {UA_SBB_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h574] = {UA_SBB_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h575] = {UA_SBB_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h576] = {UA_SBB_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h577] = {UA_SBB_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h508] = {UA_AND_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h509] = {UA_AND_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h50a] = {UA_AND_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h50b] = {UA_AND_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h50c] = {UA_AND_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h50d] = {UA_AND_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h50e] = {UA_AND_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h50f] = {UA_AND_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h510] = {UA_XOR_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h511] = {UA_XOR_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h512] = {UA_XOR_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h513] = {UA_XOR_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h514] = {UA_XOR_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h515] = {UA_XOR_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h516] = {UA_XOR_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h517] = {UA_XOR_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h518] = {UA_OR_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h519] = {UA_OR_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h51a] = {UA_OR_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h51b] = {UA_OR_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h51c] = {UA_OR_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h51d] = {UA_OR_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h51e] = {UA_OR_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h51f] = {UA_OR_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h5a0] = {UA_ADDNC_SPR_IR2_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h5a1] = {UA_ADDNC_SPR_IR2_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h5a2] = {UA_ADDNC_SPR_IR2_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h5a3] = {UA_ADDNC_SPR_IR2_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h5b0] = {UA_SUBNB_SPR_IR2_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h5b1] = {UA_SUBNB_SPR_IR2_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h5b2] = {UA_SUBNB_SPR_IR2_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h5b3] = {UA_SUBNB_SPR_IR2_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h5c0] = {UA_ADD_SPR_IR2_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h5c1] = {UA_ADD_SPR_IR2_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h5c2] = {UA_ADD_SPR_IR2_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h5c3] = {UA_ADD_SPR_IR2_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h5d0] = {UA_ADC_SPR_IR2_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h5d1] = {UA_ADC_SPR_IR2_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h5d2] = {UA_ADC_SPR_IR2_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h5d3] = {UA_ADC_SPR_IR2_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h5e0] = {UA_SUB_SPR_IR2_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h5e1] = {UA_SUB_SPR_IR2_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h5e2] = {UA_SUB_SPR_IR2_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h5e3] = {UA_SUB_SPR_IR2_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h5f0] = {UA_SBB_SPR_IR2_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h5f1] = {UA_SBB_SPR_IR2_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h5f2] = {UA_SBB_SPR_IR2_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h5f3] = {UA_SBB_SPR_IR2_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h588] = {UA_AND_SPR_IR2_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h589] = {UA_AND_SPR_IR2_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h58a] = {UA_AND_SPR_IR2_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h58b] = {UA_AND_SPR_IR2_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h590] = {UA_XOR_SPR_IR2_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h591] = {UA_XOR_SPR_IR2_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h592] = {UA_XOR_SPR_IR2_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h593] = {UA_XOR_SPR_IR2_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h598] = {UA_OR_SPR_IR2_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h599] = {UA_OR_SPR_IR2_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h59a] = {UA_OR_SPR_IR2_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h59b] = {UA_OR_SPR_IR2_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h528] = {UA_CMPBNB_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h529] = {UA_CMPBNB_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h52a] = {UA_CMPBNB_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h52b] = {UA_CMPBNB_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h52c] = {UA_CMPBNB_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h52d] = {UA_CMPBNB_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h52e] = {UA_CMPBNB_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h52f] = {UA_CMPBNB_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h538] = {UA_CMPB_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h539] = {UA_CMPB_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h53a] = {UA_CMPB_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h53b] = {UA_CMPB_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h53c] = {UA_CMPB_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h53d] = {UA_CMPB_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h53e] = {UA_CMPB_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h53f] = {UA_CMPB_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h548] = {UA_BITNZ_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h549] = {UA_BITNZ_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h54a] = {UA_BITNZ_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h54b] = {UA_BITNZ_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h54c] = {UA_BITNZ_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h54d] = {UA_BITNZ_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h54e] = {UA_BITNZ_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h54f] = {UA_BITNZ_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h558] = {UA_BITZ_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h559] = {UA_BITZ_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h55a] = {UA_BITZ_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h55b] = {UA_BITZ_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h55c] = {UA_BITZ_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h55d] = {UA_BITZ_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h55e] = {UA_BITZ_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h55f] = {UA_BITZ_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h568] = {UA_CMPNZ_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h569] = {UA_CMPNZ_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h56a] = {UA_CMPNZ_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h56b] = {UA_CMPNZ_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h56c] = {UA_CMPNZ_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h56d] = {UA_CMPNZ_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h56e] = {UA_CMPNZ_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h56f] = {UA_CMPNZ_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h578] = {UA_CMPZ_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h579] = {UA_CMPZ_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h57a] = {UA_CMPZ_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h57b] = {UA_CMPZ_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h57c] = {UA_CMPZ_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h57d] = {UA_CMPZ_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h57e] = {UA_CMPZ_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h57f] = {UA_CMPZ_RF_IR210_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h5a8] = {UA_CMPBNB_SPR_IR2_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h5a9] = {UA_CMPBNB_SPR_IR2_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h5aa] = {UA_CMPBNB_SPR_IR2_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h5ab] = {UA_CMPBNB_SPR_IR2_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h5b8] = {UA_CMPB_SPR_IR2_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h5b9] = {UA_CMPB_SPR_IR2_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h5ba] = {UA_CMPB_SPR_IR2_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h5bb] = {UA_CMPB_SPR_IR2_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h5c8] = {UA_BITNZ_SPR_IR2_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h5c9] = {UA_BITNZ_SPR_IR2_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h5ca] = {UA_BITNZ_SPR_IR2_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h5cb] = {UA_BITNZ_SPR_IR2_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h5d8] = {UA_BITZ_SPR_IR2_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h5d9] = {UA_BITZ_SPR_IR2_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h5da] = {UA_BITZ_SPR_IR2_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h5db] = {UA_BITZ_SPR_IR2_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h5e8] = {UA_CMPNZ_SPR_IR2_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h5e9] = {UA_CMPNZ_SPR_IR2_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h5ea] = {UA_CMPNZ_SPR_IR2_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h5eb] = {UA_CMPNZ_SPR_IR2_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h5f8] = {UA_CMPZ_SPR_IR2_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h5f9] = {UA_CMPZ_SPR_IR2_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h5fa] = {UA_CMPZ_SPR_IR2_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h5fb] = {UA_CMPZ_SPR_IR2_IMM, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h668] = {UA_LD_IR210_ABS, 1'd0, 2'd2, ISEFM_NONE};
    ird_lut['h669] = {UA_LD_IR210_ABS, 1'd0, 2'd2, ISEFM_NONE};
    ird_lut['h66a] = {UA_LD_IR210_ABS, 1'd0, 2'd2, ISEFM_NONE};
    ird_lut['h66b] = {UA_LD_IR210_ABS, 1'd0, 2'd2, ISEFM_NONE};
    ird_lut['h66c] = {UA_LD_IR210_ABS, 1'd0, 2'd2, ISEFM_NONE};
    ird_lut['h66d] = {UA_LD_IR210_ABS, 1'd0, 2'd2, ISEFM_NONE};
    ird_lut['h66e] = {UA_LD_IR210_ABS, 1'd0, 2'd2, ISEFM_NONE};
    ird_lut['h66f] = {UA_LD_IR210_ABS, 1'd0, 2'd2, ISEFM_NONE};
    ird_lut['h60f] = {UA_LSPD, 1'd0, 2'd2, ISEFM_NONE};
    ird_lut['h61f] = {UA_LBCD, 1'd0, 2'd2, ISEFM_NONE};
    ird_lut['h62f] = {UA_LDED, 1'd0, 2'd2, ISEFM_NONE};
    ird_lut['h63f] = {UA_LHLD, 1'd0, 2'd2, ISEFM_NONE};
    ird_lut['h678] = {UA_ST_IR210_ABS, 1'd0, 2'd2, ISEFM_NONE};
    ird_lut['h679] = {UA_ST_IR210_ABS, 1'd0, 2'd2, ISEFM_NONE};
    ird_lut['h67a] = {UA_ST_IR210_ABS, 1'd0, 2'd2, ISEFM_NONE};
    ird_lut['h67b] = {UA_ST_IR210_ABS, 1'd0, 2'd2, ISEFM_NONE};
    ird_lut['h67c] = {UA_ST_IR210_ABS, 1'd0, 2'd2, ISEFM_NONE};
    ird_lut['h67d] = {UA_ST_IR210_ABS, 1'd0, 2'd2, ISEFM_NONE};
    ird_lut['h67e] = {UA_ST_IR210_ABS, 1'd0, 2'd2, ISEFM_NONE};
    ird_lut['h67f] = {UA_ST_IR210_ABS, 1'd0, 2'd2, ISEFM_NONE};
    ird_lut['h60e] = {UA_SSPD, 1'd0, 2'd2, ISEFM_NONE};
    ird_lut['h61e] = {UA_SBCD, 1'd0, 2'd2, ISEFM_NONE};
    ird_lut['h62e] = {UA_SDED, 1'd0, 2'd2, ISEFM_NONE};
    ird_lut['h63e] = {UA_SHLD, 1'd0, 2'd2, ISEFM_NONE};
    ird_lut['h6a1] = {UA_ADDNC_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6a2] = {UA_ADDNC_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6a3] = {UA_ADDNC_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6a4] = {UA_ADDNC_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6a5] = {UA_ADDNC_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6a6] = {UA_ADDNC_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6a7] = {UA_ADDNC_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6b1] = {UA_SUBNB_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6b2] = {UA_SUBNB_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6b3] = {UA_SUBNB_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6b4] = {UA_SUBNB_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6b5] = {UA_SUBNB_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6b6] = {UA_SUBNB_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6b7] = {UA_SUBNB_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6c1] = {UA_ADD_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6c2] = {UA_ADD_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6c3] = {UA_ADD_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6c4] = {UA_ADD_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6c5] = {UA_ADD_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6c6] = {UA_ADD_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6c7] = {UA_ADD_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6d1] = {UA_ADC_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6d2] = {UA_ADC_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6d3] = {UA_ADC_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6d4] = {UA_ADC_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6d5] = {UA_ADC_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6d6] = {UA_ADC_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6d7] = {UA_ADC_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6e1] = {UA_SUB_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6e2] = {UA_SUB_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6e3] = {UA_SUB_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6e4] = {UA_SUB_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6e5] = {UA_SUB_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6e6] = {UA_SUB_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6e7] = {UA_SUB_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6f1] = {UA_SBB_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6f2] = {UA_SBB_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6f3] = {UA_SBB_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6f4] = {UA_SBB_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6f5] = {UA_SBB_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6f6] = {UA_SBB_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6f7] = {UA_SBB_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h689] = {UA_AND_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h68a] = {UA_AND_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h68b] = {UA_AND_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h68c] = {UA_AND_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h68d] = {UA_AND_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h68e] = {UA_AND_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h68f] = {UA_AND_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h691] = {UA_XOR_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h692] = {UA_XOR_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h693] = {UA_XOR_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h694] = {UA_XOR_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h695] = {UA_XOR_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h696] = {UA_XOR_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h697] = {UA_XOR_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h699] = {UA_OR_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h69a] = {UA_OR_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h69b] = {UA_OR_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h69c] = {UA_OR_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h69d] = {UA_OR_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h69e] = {UA_OR_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h69f] = {UA_OR_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6a9] = {UA_CMPBNB_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6aa] = {UA_CMPBNB_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6ab] = {UA_CMPBNB_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6ac] = {UA_CMPBNB_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6ad] = {UA_CMPBNB_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6ae] = {UA_CMPBNB_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6af] = {UA_CMPBNB_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6b9] = {UA_CMPB_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6ba] = {UA_CMPB_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6bb] = {UA_CMPB_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6bc] = {UA_CMPB_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6bd] = {UA_CMPB_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6be] = {UA_CMPB_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6bf] = {UA_CMPB_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6c9] = {UA_BITNZ_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6ca] = {UA_BITNZ_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6cb] = {UA_BITNZ_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6cc] = {UA_BITNZ_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6cd] = {UA_BITNZ_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6ce] = {UA_BITNZ_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6cf] = {UA_BITNZ_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6d9] = {UA_BITZ_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6da] = {UA_BITZ_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6db] = {UA_BITZ_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6dc] = {UA_BITZ_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6dd] = {UA_BITZ_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6de] = {UA_BITZ_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6df] = {UA_BITZ_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6e9] = {UA_CMPNZ_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6ea] = {UA_CMPNZ_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6eb] = {UA_CMPNZ_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6ec] = {UA_CMPNZ_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6ed] = {UA_CMPNZ_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6ee] = {UA_CMPNZ_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6ef] = {UA_CMPNZ_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6f9] = {UA_CMPZ_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6fa] = {UA_CMPZ_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6fb] = {UA_CMPZ_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6fc] = {UA_CMPZ_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6fd] = {UA_CMPZ_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6fe] = {UA_CMPZ_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h6ff] = {UA_CMPZ_A_IND, 1'd0, 2'd0, ISEFM_NONE};
    ird_lut['h7a0] = {UA_ADDNC_A_WA, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h7b0] = {UA_SUBNB_A_WA, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h7c0] = {UA_ADD_A_WA, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h7d0] = {UA_ADC_A_WA, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h7e0] = {UA_SUB_A_WA, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h7f0] = {UA_SBB_A_WA, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h788] = {UA_AND_A_WA, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h790] = {UA_XOR_A_WA, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h798] = {UA_OR_A_WA, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h7a8] = {UA_CMPBNB_A_WA, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h7b8] = {UA_CMPB_A_WA, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h7c8] = {UA_BITNZ_A_WA, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h7d8] = {UA_BITZ_A_WA, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h7e8] = {UA_CMPNZ_A_WA, 1'd0, 2'd1, ISEFM_NONE};
    ird_lut['h7f8] = {UA_CMPZ_A_WA, 1'd0, 2'd1, ISEFM_NONE};
