typedef enum reg [9:0]
{
    UA_IDLE,
    UA_SKIP_OP2,
    UA__2,
    UA__3,
    UA_SKIP_OP1,
    UA__5,
    UA__6,
    UA_MOV_A_RF_IR210,
    UA__8,
    UA__9,
    UA_MOV_RF_IR210_A,
    UA__B,
    UA__C,
    UA_MOV_RF_IR210_IMM,
    UA__E,
    UA__F,
    UA_LD_A_WA,
    UA__11,
    UA__12,
    UA__13,
    UA__14,
    UA__15,
    UA_LDX_SP_IMM,
    UA__17,
    UA__18,
    UA__19,
    UA__1A,
    UA__1B,
    UA_LDX_BC_IMM,
    UA__1D,
    UA__1E,
    UA__1F,
    UA__20,
    UA__21,
    UA_LDX_DE_IMM,
    UA__23,
    UA__24,
    UA__25,
    UA__26,
    UA__27,
    UA_LDX_HL_IMM,
    UA__29,
    UA__2A,
    UA__2B,
    UA__2C,
    UA__2D,
    UA_LDAX,
    UA__2F,
    UA__30,
    UA_STX_A,
    UA__32,
    UA__33,
    UA_STX_RF_W,
    UA__35,
    UA__36,
    UA__37,
    UA__38,
    UA__39,
    UA_STW_A,
    UA__3B,
    UA__3C,
    UA__3D,
    UA__3E,
    UA__3F,
    UA_STW_IMM,
    UA__41,
    UA__42,
    UA__43,
    UA__44,
    UA__45,
    UA__46,
    UA__47,
    UA__48,
    UA_TABLE,
    UA__4A,
    UA__4B,
    UA__4C,
    UA__4D,
    UA__4E,
    UA__4F,
    UA__50,
    UA__51,
    UA__52,
    UA__53,
    UA__54,
    UA__55,
    UA__56,
    UA__57,
    UA_BLOCK,
    UA__59,
    UA__5A,
    UA__5B,
    UA__5C,
    UA__5D,
    UA__5E,
    UA__5F,
    UA__60,
    UA_AND_WA_IMM,
    UA__62,
    UA__63,
    UA__64,
    UA__65,
    UA__66,
    UA__67,
    UA__68,
    UA__69,
    UA__6A,
    UA__6B,
    UA__6C,
    UA_OR_WA_IMM,
    UA__6E,
    UA__6F,
    UA__70,
    UA__71,
    UA__72,
    UA__73,
    UA__74,
    UA__75,
    UA__76,
    UA__77,
    UA__78,
    UA_AND_A_IMM,
    UA__7A,
    UA__7B,
    UA__7C,
    UA_XOR_A_IMM,
    UA__7E,
    UA__7F,
    UA__80,
    UA_OR_A_IMM,
    UA__82,
    UA__83,
    UA__84,
    UA_ON_WA_IMM,
    UA__86,
    UA__87,
    UA__88,
    UA__89,
    UA__8A,
    UA__8B,
    UA__8C,
    UA__8D,
    UA__8E,
    UA_NEQ_WA_IMM,
    UA__90,
    UA__91,
    UA__92,
    UA__93,
    UA__94,
    UA__95,
    UA__96,
    UA__97,
    UA__98,
    UA_GT_A_IMM,
    UA__9A,
    UA__9B,
    UA__9C,
    UA_LT_A_IMM,
    UA__9E,
    UA__9F,
    UA__A0,
    UA_ON_A_IMM,
    UA__A2,
    UA__A3,
    UA__A4,
    UA_OFF_A_IMM,
    UA__A6,
    UA__A7,
    UA__A8,
    UA_NEQ_A_IMM,
    UA__AA,
    UA__AB,
    UA__AC,
    UA_EQ_A_IMM,
    UA__AE,
    UA__AF,
    UA__B0,
    UA_ADDNC_A_IMM,
    UA__B2,
    UA__B3,
    UA__B4,
    UA_SUBNB_A_IMM,
    UA__B6,
    UA__B7,
    UA__B8,
    UA_ADD_A_IMM,
    UA__BA,
    UA__BB,
    UA__BC,
    UA_ADC_A_IMM,
    UA__BE,
    UA__BF,
    UA__C0,
    UA_SUB_A_IMM,
    UA__C2,
    UA__C3,
    UA__C4,
    UA_SBB_A_IMM,
    UA__C6,
    UA__C7,
    UA__C8,
    UA_INCR_WA,
    UA__CA,
    UA__CB,
    UA__CC,
    UA__CD,
    UA__CE,
    UA__CF,
    UA__D0,
    UA__D1,
    UA_DECR_WA,
    UA__D3,
    UA__D4,
    UA__D5,
    UA__D6,
    UA__D7,
    UA__D8,
    UA__D9,
    UA__DA,
    UA_INCR_RF_IR210,
    UA__DC,
    UA_DECR_RF_IR210,
    UA__DE,
    UA_INC_SP,
    UA__E0,
    UA__E1,
    UA_INC_BC,
    UA__E3,
    UA__E4,
    UA_INC_DE,
    UA__E6,
    UA__E7,
    UA_INC_HL,
    UA__E9,
    UA__EA,
    UA_DEC_SP,
    UA__EC,
    UA__ED,
    UA_DEC_BC,
    UA__EF,
    UA__F0,
    UA_DEC_DE,
    UA__F2,
    UA__F3,
    UA_DEC_HL,
    UA__F5,
    UA__F6,
    UA_DAA,
    UA__F8,
    UA_JR,
    UA__FA,
    UA__FB,
    UA__FC,
    UA__FD,
    UA__FE,
    UA__FF,
    UA__100,
    UA__101,
    UA_JRE_P,
    UA__103,
    UA__104,
    UA__105,
    UA__106,
    UA__107,
    UA__108,
    UA__109,
    UA__10A,
    UA_JRE_N,
    UA__10C,
    UA__10D,
    UA__10E,
    UA__10F,
    UA__110,
    UA__111,
    UA__112,
    UA__113,
    UA_JMP,
    UA__115,
    UA__116,
    UA__117,
    UA__118,
    UA__119,
    UA_JB,
    UA_CALF,
    UA__11C,
    UA__11D,
    UA__11E,
    UA__11F,
    UA__120,
    UA__121,
    UA__122,
    UA__123,
    UA__124,
    UA__125,
    UA__126,
    UA_CALT,
    UA__128,
    UA__129,
    UA__12A,
    UA__12B,
    UA__12C,
    UA__12D,
    UA__12E,
    UA__12F,
    UA__130,
    UA__131,
    UA__132,
    UA__133,
    UA__134,
    UA__135,
    UA_INT,
    UA__137,
    UA__138,
    UA__139,
    UA__13A,
    UA__13B,
    UA__13C,
    UA__13D,
    UA__13E,
    UA__13F,
    UA__140,
    UA__141,
    UA__142,
    UA__143,
    UA__144,
    UA__145,
    UA__146,
    UA__147,
    UA_RET,
    UA__149,
    UA__14A,
    UA__14B,
    UA__14C,
    UA__14D,
    UA_RETI,
    UA__14F,
    UA__150,
    UA__151,
    UA__152,
    UA__153,
    UA__154,
    UA__155,
    UA__156,
    UA_BIT,
    UA__158,
    UA__159,
    UA__15A,
    UA__15B,
    UA__15C,
    UA__15D,
    UA_STM,
    UA_RLL_A_,
    UA__160,
    UA__161,
    UA_RLR_A_,
    UA__163,
    UA__164,
    UA_RLL_C_,
    UA__166,
    UA__167,
    UA_RLR_C_,
    UA__169,
    UA__16A,
    UA_SLL_A_,
    UA__16C,
    UA__16D,
    UA_SLR_A_,
    UA__16F,
    UA__170,
    UA_SLL_C_,
    UA__172,
    UA__173,
    UA_SLR_C_,
    UA__175,
    UA__176,
    UA_PUSH_VA,
    UA__178,
    UA__179,
    UA__17A,
    UA__17B,
    UA__17C,
    UA__17D,
    UA__17E,
    UA__17F,
    UA_POP_VA,
    UA__181,
    UA__182,
    UA__183,
    UA__184,
    UA__185,
    UA_PUSH_BC,
    UA__187,
    UA__188,
    UA__189,
    UA__18A,
    UA__18B,
    UA__18C,
    UA__18D,
    UA__18E,
    UA_POP_BC,
    UA__190,
    UA__191,
    UA__192,
    UA__193,
    UA__194,
    UA_PUSH_DE,
    UA__196,
    UA__197,
    UA__198,
    UA__199,
    UA__19A,
    UA__19B,
    UA__19C,
    UA__19D,
    UA_POP_DE,
    UA__19F,
    UA__1A0,
    UA__1A1,
    UA__1A2,
    UA__1A3,
    UA_PUSH_HL,
    UA__1A5,
    UA__1A6,
    UA__1A7,
    UA__1A8,
    UA__1A9,
    UA__1AA,
    UA__1AB,
    UA__1AC,
    UA_POP_HL,
    UA__1AE,
    UA__1AF,
    UA__1B0,
    UA__1B1,
    UA__1B2,
    UA_SKIP_I,
    UA_SKIP_C,
    UA_SKIP_NI,
    UA_SKIP_NC,
    UA_EI,
    UA_DI,
    UA_MOV_A_SPR_IR3,
    UA__1BA,
    UA__1BB,
    UA_MOV_SPR_IR3_A,
    UA__1BD,
    UA__1BE,
    UA_ADDNC_RF_IR210_A,
    UA__1C0,
    UA__1C1,
    UA_SUBNB_RF_IR210_A,
    UA__1C3,
    UA__1C4,
    UA_ADD_RF_IR210_A,
    UA__1C6,
    UA__1C7,
    UA_ADC_RF_IR210_A,
    UA__1C9,
    UA__1CA,
    UA_SUB_RF_IR210_A,
    UA__1CC,
    UA__1CD,
    UA_SBB_RF_IR210_A,
    UA__1CF,
    UA__1D0,
    UA_ADDNC_A_RF_IR210,
    UA__1D2,
    UA__1D3,
    UA_SUBNB_A_RF_IR210,
    UA__1D5,
    UA__1D6,
    UA_ADD_A_RF_IR210,
    UA__1D8,
    UA__1D9,
    UA_ADC_A_RF_IR210,
    UA__1DB,
    UA__1DC,
    UA_SUB_A_RF_IR210,
    UA__1DE,
    UA__1DF,
    UA_SBB_A_RF_IR210,
    UA__1E1,
    UA__1E2,
    UA_ADDNC_RF_IR210_IMM,
    UA__1E4,
    UA__1E5,
    UA__1E6,
    UA_SUBNB_RF_IR210_IMM,
    UA__1E8,
    UA__1E9,
    UA__1EA,
    UA_ADD_RF_IR210_IMM,
    UA__1EC,
    UA__1ED,
    UA__1EE,
    UA_ADC_RF_IR210_IMM,
    UA__1F0,
    UA__1F1,
    UA__1F2,
    UA_OFF_RF_IR210_IMM,
    UA__1F4,
    UA__1F5,
    UA__1F6,
    UA_SUB_RF_IR210_IMM,
    UA__1F8,
    UA__1F9,
    UA__1FA,
    UA_SBB_RF_IR210_IMM,
    UA__1FC,
    UA__1FD,
    UA__1FE,
    UA_AND_SPR_IR2_IMM,
    UA__200,
    UA__201,
    UA__202,
    UA_XOR_SPR_IR2_IMM,
    UA__204,
    UA__205,
    UA__206,
    UA_OR_SPR_IR2_IMM,
    UA__208,
    UA__209,
    UA__20A,
    UA_ON_RF_IR210_IMM,
    UA__20C,
    UA__20D,
    UA__20E,
    UA_ON_SPR_IR2_IMM,
    UA__210,
    UA__211,
    UA__212,
    UA_OFF_SPR_IR2_IMM,
    UA__214,
    UA__215,
    UA__216,
    UA_LD_IR210_ABS,
    UA__218,
    UA__219,
    UA__21A,
    UA__21B,
    UA__21C,
    UA__21D,
    UA__21E,
    UA__21F,
    UA_ST_IR210_ABS,
    UA__221,
    UA__222,
    UA__223,
    UA__224,
    UA__225,
    UA__226,
    UA__227,
    UA__228,
    UA_ADD,
    UA__22A,
    UA__22B,
    UA__22C,
    UA_SUB,
    UA__22E,
    UA__22F,
    UA__230,
    UA_ADD_A_WA,
    UA__232,
    UA__233,
    UA__234,
    UA__235,
    UA__236,
    UA__237,
    UA_AND_A_WA,
    UA__239,
    UA__23A,
    UA__23B,
    UA__23C,
    UA__23D,
    UA__23E,
    UA_OR_A_WA,
    UA__240,
    UA__241,
    UA__242,
    UA__243,
    UA__244,
    UA__245
} e_uaddr;    // ucode address

typedef reg [7:0] t_naddr;    // ncode address

typedef enum reg [1:0]
{
    UBM_ADV,
    UBM_END,
    UBM_DA
} e_ubm;    // branch mode

typedef enum reg [1:0]
{
    UTX_T1,
    UTX_T2,
    UTX_T3,
    UTX_T4
} e_mcy;    // machine cycle

typedef enum reg [3:0]
{
    URFS_V,
    URFS_A,
    URFS_B,
    URFS_C,
    URFS_D,
    URFS_E,
    URFS_H,
    URFS_L,
    URFS_PSW,
    URFS_SPL,
    URFS_SPH,
    URFS_PCL,
    URFS_PCH,
    URFS_IR210,
    URFS_W
} e_urfs;    // register file select

typedef enum reg [2:0]
{
    UIDBS_0,
    UIDBS_RF,
    UIDBS_DB,
    UIDBS_CO,
    UIDBS_SPR,
    UIDBS_SDG
} e_idbs;    // idb select

typedef enum reg [3:0]
{
    ULTS_NONE,
    ULTS_RF,
    ULTS_DOR,
    ULTS_AI,
    ULTS_BI,
    ULTS_IE,
    ULTS_SPR
} e_lts;    // load target select

typedef enum reg [3:0]
{
    UABS_PC,
    UABS_SP,
    UABS_BC,
    UABS_DE,
    UABS_HL,
    UABS_VW,
    UABS_IDB_W,
    UABS_IR210,
    UABS_AOR,
    UABS_NABI
} e_abs;    // ab select

typedef enum reg [3:0]
{
    USPR_PA,
    USPR_PB,
    USPR_PC,
    USPR_MK,
    USPR_MB,
    USPR_MC,
    USPR_TM0,
    USPR_TM1,
    USPR_S,
    USPR_TMM
} e_spr;    // special register

typedef enum reg [0:0]
{
    USRS_IR2,
    USRS_IR3
} e_sprs;    // special register select

typedef enum reg [2:0]
{
    USDGS_JRL,
    USDGS_JRH,
    USDGS_CALF,
    USDGS_CALT,
    USDGS_INTVA,
    USDGS_BIT
} e_sdgs;    // special data generator select

typedef enum reg [3:0]
{
    UAO_NOP,
    UAO_SUM,
    UAO_INC,
    UAO_DEC,
    UAO_OR,
    UAO_AND,
    UAO_EOR,
    UAO_LSL,
    UAO_ROL,
    UAO_LSR,
    UAO_ROR
} e_aluop;    // ALU operation

typedef enum reg [1:0]
{
    UCIS_0,
    UCIS_1,
    UCIS_CCO,
    UCIS_PSW_CY
} e_cis;    // ALU carry in select

typedef enum reg [3:0]
{
    USKS_PSW_SK,
    USKS_1,
    USKS_C,
    USKS_NC,
    USKS_Z,
    USKS_NZ,
    USKS_I,
    USKS_NI,
    USKS_0
} e_sks;    // SKip flag source

typedef struct packed
{
    e_uaddr uaddr;    // microcode entry point
    reg [0:0] m1_overlap;    // New M1 starts immediately
    reg [1:0] skipn;    // Number of operands to skip when ins. is skipped
} s_ird;

typedef struct packed
{
    t_naddr naddr;    // nanocode address
    e_ubm bm;    // branch mode
    reg [0:0] m1;    // Fetch next opcode (start M1)
} s_uc;

typedef struct packed
{
    reg [2:0] idx;    // general-purpose data
    e_urfs rfos;    // register file output select -> idb
    e_urfs rfts;    // register file target select
    e_idbs idbs;    // idb select
    e_lts lts;    // load target select
    e_abs abs;    // ab select
    e_abs abits;    // abi target select
    reg [0:0] pc_inc;    // increment PC
    reg [0:0] ab_inc;    // increment ab
    reg [0:0] ab_dec;    // decrement ab
    reg [0:0] aout;    // ab -> AOR
    reg [0:0] load;    // assert RDB (read operation)
    reg [0:0] store;    // dor -> DB
    e_aluop aluop;    // ALU operation
    e_cis cis;    // ALU carry in select
    reg [0:0] bi0;    // Zero BI
    reg [0:0] bin;    // Negate BI
    reg [0:0] pswz;    // (CO == 0) -> PSW.Z
    reg [0:0] pswcy;    // CCO -> PSW.CY
    reg [0:0] pswhc;    // CHO -> PSW.HC
    e_sks pswsk;    // PSW.SK source
    e_sprs sprs;    // special register select
    e_sdgs sdgs;    // special data generator select
    reg [0:0] daa;    // decimal adjust const -> BI
    reg [0:0] rpir;    // IR[2:0] selects reg. pair and inc/dec
} s_nc;

