s_uc urom [1030];
initial begin
  urom[   0] = 10'b0000000010;
  urom[   1] = 10'b0000000100;
  urom[   2] = 10'b0000001000;
  urom[   3] = 10'b0000000000;
  urom[   4] = 10'b0000000100;
  urom[   5] = 10'b0000001000;
  urom[   6] = 10'b0000000011;
  urom[   7] = 10'b0000010000;
  urom[   8] = 10'b0000000000;
  urom[   9] = 10'b0000010110;
  urom[  10] = 10'b0000011000;
  urom[  11] = 10'b0000000000;
  urom[  12] = 10'b0000010110;
  urom[  13] = 10'b0000000100;
  urom[  14] = 10'b0000001000;
  urom[  15] = 10'b0000011111;
  urom[  16] = 10'b0000000100;
  urom[  17] = 10'b0000001000;
  urom[  18] = 10'b0000011111;
  urom[  19] = 10'b0000000100;
  urom[  20] = 10'b0000001000;
  urom[  21] = 10'b0000011111;
  urom[  22] = 10'b0000000100;
  urom[  23] = 10'b0000001000;
  urom[  24] = 10'b0000100000;
  urom[  25] = 10'b0000100100;
  urom[  26] = 10'b0000001000;
  urom[  27] = 10'b0000101011;
  urom[  28] = 10'b0000000100;
  urom[  29] = 10'b0000001000;
  urom[  30] = 10'b0000101100;
  urom[  31] = 10'b0000000100;
  urom[  32] = 10'b0000001000;
  urom[  33] = 10'b0000110011;
  urom[  34] = 10'b0000000100;
  urom[  35] = 10'b0000001000;
  urom[  36] = 10'b0000110100;
  urom[  37] = 10'b0000000100;
  urom[  38] = 10'b0000001000;
  urom[  39] = 10'b0000111011;
  urom[  40] = 10'b0000000100;
  urom[  41] = 10'b0000001000;
  urom[  42] = 10'b0000111100;
  urom[  43] = 10'b0000000100;
  urom[  44] = 10'b0000001000;
  urom[  45] = 10'b0001000011;
  urom[  46] = 10'b0000000100;
  urom[  47] = 10'b0000001000;
  urom[  48] = 10'b0001000100;
  urom[  49] = 10'b0000000100;
  urom[  50] = 10'b0000001000;
  urom[  51] = 10'b0001001011;
  urom[  52] = 10'b0001001100;
  urom[  53] = 10'b0000001000;
  urom[  54] = 10'b0000101011;
  urom[  55] = 10'b0001010000;
  urom[  56] = 10'b0000001100;
  urom[  57] = 10'b0000010111;
  urom[  58] = 10'b0000000100;
  urom[  59] = 10'b0000001000;
  urom[  60] = 10'b0000100000;
  urom[  61] = 10'b0001010100;
  urom[  62] = 10'b0000001100;
  urom[  63] = 10'b0000010111;
  urom[  64] = 10'b0000000100;
  urom[  65] = 10'b0000001000;
  urom[  66] = 10'b0000100000;
  urom[  67] = 10'b0001011000;
  urom[  68] = 10'b0000001100;
  urom[  69] = 10'b0000010111;
  urom[  70] = 10'b0000000100;
  urom[  71] = 10'b0000001000;
  urom[  72] = 10'b0000100000;
  urom[  73] = 10'b0000000100;
  urom[  74] = 10'b0000001000;
  urom[  75] = 10'b0001011100;
  urom[  76] = 10'b0001100000;
  urom[  77] = 10'b0000001100;
  urom[  78] = 10'b0000010111;
  urom[  79] = 10'b0001100100;
  urom[  80] = 10'b0000000000;
  urom[  81] = 10'b0000000000;
  urom[  82] = 10'b0001101000;
  urom[  83] = 10'b0001101100;
  urom[  84] = 10'b0000000000;
  urom[  85] = 10'b0001110000;
  urom[  86] = 10'b0000000000;
  urom[  87] = 10'b0000000000;
  urom[  88] = 10'b0001110100;
  urom[  89] = 10'b0000001000;
  urom[  90] = 10'b0001111000;
  urom[  91] = 10'b0001111100;
  urom[  92] = 10'b0000001000;
  urom[  93] = 10'b0000111011;
  urom[  94] = 10'b0010000000;
  urom[  95] = 10'b0010000100;
  urom[  96] = 10'b0000100000;
  urom[  97] = 10'b0010001000;
  urom[  98] = 10'b0010001100;
  urom[  99] = 10'b0000000000;
  urom[ 100] = 10'b0010010000;
  urom[ 101] = 10'b0010010100;
  urom[ 102] = 10'b0010011011;
  urom[ 103] = 10'b0010011110;
  urom[ 104] = 10'b0010100010;
  urom[ 105] = 10'b0000000100;
  urom[ 106] = 10'b0000001000;
  urom[ 107] = 10'b0000100000;
  urom[ 108] = 10'b0000100100;
  urom[ 109] = 10'b0000001000;
  urom[ 110] = 10'b0010100100;
  urom[ 111] = 10'b0000000100;
  urom[ 112] = 10'b0000001000;
  urom[ 113] = 10'b0010101000;
  urom[ 114] = 10'b0001100000;
  urom[ 115] = 10'b0000001100;
  urom[ 116] = 10'b0010101111;
  urom[ 117] = 10'b0000000100;
  urom[ 118] = 10'b0000001000;
  urom[ 119] = 10'b0000100000;
  urom[ 120] = 10'b0000100100;
  urom[ 121] = 10'b0000001000;
  urom[ 122] = 10'b0010100100;
  urom[ 123] = 10'b0000000100;
  urom[ 124] = 10'b0000001000;
  urom[ 125] = 10'b0010110000;
  urom[ 126] = 10'b0001100000;
  urom[ 127] = 10'b0000001100;
  urom[ 128] = 10'b0010101111;
  urom[ 129] = 10'b0010110100;
  urom[ 130] = 10'b0000001000;
  urom[ 131] = 10'b0010101001;
  urom[ 132] = 10'b0010111010;
  urom[ 133] = 10'b0010110100;
  urom[ 134] = 10'b0000001000;
  urom[ 135] = 10'b0010111101;
  urom[ 136] = 10'b0010111010;
  urom[ 137] = 10'b0010110100;
  urom[ 138] = 10'b0000001000;
  urom[ 139] = 10'b0010110001;
  urom[ 140] = 10'b0010111010;
  urom[ 141] = 10'b0000000100;
  urom[ 142] = 10'b0000001000;
  urom[ 143] = 10'b0000100000;
  urom[ 144] = 10'b0000100100;
  urom[ 145] = 10'b0000001000;
  urom[ 146] = 10'b0010100100;
  urom[ 147] = 10'b0000000100;
  urom[ 148] = 10'b0000001000;
  urom[ 149] = 10'b0011000001;
  urom[ 150] = 10'b0011000110;
  urom[ 151] = 10'b0000000100;
  urom[ 152] = 10'b0000001000;
  urom[ 153] = 10'b0000100000;
  urom[ 154] = 10'b0000100100;
  urom[ 155] = 10'b0000001000;
  urom[ 156] = 10'b0010100100;
  urom[ 157] = 10'b0000000100;
  urom[ 158] = 10'b0000001000;
  urom[ 159] = 10'b0011001001;
  urom[ 160] = 10'b0011001110;
  urom[ 161] = 10'b0000000100;
  urom[ 162] = 10'b0000001000;
  urom[ 163] = 10'b0000100000;
  urom[ 164] = 10'b0000100100;
  urom[ 165] = 10'b0000001000;
  urom[ 166] = 10'b0010100100;
  urom[ 167] = 10'b0000000100;
  urom[ 168] = 10'b0000001000;
  urom[ 169] = 10'b0010101001;
  urom[ 170] = 10'b0011010010;
  urom[ 171] = 10'b0000000100;
  urom[ 172] = 10'b0000001000;
  urom[ 173] = 10'b0000100000;
  urom[ 174] = 10'b0000100100;
  urom[ 175] = 10'b0000001000;
  urom[ 176] = 10'b0010100100;
  urom[ 177] = 10'b0000000100;
  urom[ 178] = 10'b0000001000;
  urom[ 179] = 10'b0010101001;
  urom[ 180] = 10'b0011010110;
  urom[ 181] = 10'b0000000100;
  urom[ 182] = 10'b0000001000;
  urom[ 183] = 10'b0000100000;
  urom[ 184] = 10'b0000100100;
  urom[ 185] = 10'b0000001000;
  urom[ 186] = 10'b0010100100;
  urom[ 187] = 10'b0000000100;
  urom[ 188] = 10'b0000001000;
  urom[ 189] = 10'b0011001001;
  urom[ 190] = 10'b0011011010;
  urom[ 191] = 10'b0000000100;
  urom[ 192] = 10'b0000001000;
  urom[ 193] = 10'b0000100000;
  urom[ 194] = 10'b0000100100;
  urom[ 195] = 10'b0000001000;
  urom[ 196] = 10'b0010100100;
  urom[ 197] = 10'b0000000100;
  urom[ 198] = 10'b0000001000;
  urom[ 199] = 10'b0011001001;
  urom[ 200] = 10'b0011011110;
  urom[ 201] = 10'b0010110100;
  urom[ 202] = 10'b0000001000;
  urom[ 203] = 10'b0011000001;
  urom[ 204] = 10'b0011000110;
  urom[ 205] = 10'b0010110100;
  urom[ 206] = 10'b0000001000;
  urom[ 207] = 10'b0011001001;
  urom[ 208] = 10'b0011001110;
  urom[ 209] = 10'b0010110100;
  urom[ 210] = 10'b0000001000;
  urom[ 211] = 10'b0010101001;
  urom[ 212] = 10'b0011010010;
  urom[ 213] = 10'b0010110100;
  urom[ 214] = 10'b0000001000;
  urom[ 215] = 10'b0010101001;
  urom[ 216] = 10'b0011010110;
  urom[ 217] = 10'b0010110100;
  urom[ 218] = 10'b0000001000;
  urom[ 219] = 10'b0011001001;
  urom[ 220] = 10'b0011011010;
  urom[ 221] = 10'b0010110100;
  urom[ 222] = 10'b0000001000;
  urom[ 223] = 10'b0011001001;
  urom[ 224] = 10'b0011011110;
  urom[ 225] = 10'b0010110100;
  urom[ 226] = 10'b0000001000;
  urom[ 227] = 10'b0011100001;
  urom[ 228] = 10'b0011100110;
  urom[ 229] = 10'b0010110100;
  urom[ 230] = 10'b0000001000;
  urom[ 231] = 10'b0011101001;
  urom[ 232] = 10'b0011100110;
  urom[ 233] = 10'b0010110100;
  urom[ 234] = 10'b0000001000;
  urom[ 235] = 10'b0011100001;
  urom[ 236] = 10'b0011101110;
  urom[ 237] = 10'b0010110100;
  urom[ 238] = 10'b0000001000;
  urom[ 239] = 10'b0011110001;
  urom[ 240] = 10'b0011101110;
  urom[ 241] = 10'b0010110100;
  urom[ 242] = 10'b0000001000;
  urom[ 243] = 10'b0011101001;
  urom[ 244] = 10'b0011101110;
  urom[ 245] = 10'b0010110100;
  urom[ 246] = 10'b0000001000;
  urom[ 247] = 10'b0011110101;
  urom[ 248] = 10'b0011101110;
  urom[ 249] = 10'b0000000100;
  urom[ 250] = 10'b0000001000;
  urom[ 251] = 10'b0000100000;
  urom[ 252] = 10'b0000100100;
  urom[ 253] = 10'b0000001000;
  urom[ 254] = 10'b0011111000;
  urom[ 255] = 10'b0001100000;
  urom[ 256] = 10'b0000001100;
  urom[ 257] = 10'b0011111111;
  urom[ 258] = 10'b0000000100;
  urom[ 259] = 10'b0000001000;
  urom[ 260] = 10'b0000100000;
  urom[ 261] = 10'b0000100100;
  urom[ 262] = 10'b0000001000;
  urom[ 263] = 10'b0100000000;
  urom[ 264] = 10'b0001100000;
  urom[ 265] = 10'b0000001100;
  urom[ 266] = 10'b0011111111;
  urom[ 267] = 10'b0100000100;
  urom[ 268] = 10'b0100001010;
  urom[ 269] = 10'b0100001100;
  urom[ 270] = 10'b0100001010;
  urom[ 271] = 10'b0100010000;
  urom[ 272] = 10'b0000000000;
  urom[ 273] = 10'b0000010111;
  urom[ 274] = 10'b0100010100;
  urom[ 275] = 10'b0000000000;
  urom[ 276] = 10'b0000010111;
  urom[ 277] = 10'b0100011000;
  urom[ 278] = 10'b0000000000;
  urom[ 279] = 10'b0000010111;
  urom[ 280] = 10'b0100011100;
  urom[ 281] = 10'b0000000000;
  urom[ 282] = 10'b0000010111;
  urom[ 283] = 10'b0100100000;
  urom[ 284] = 10'b0000000000;
  urom[ 285] = 10'b0000010111;
  urom[ 286] = 10'b0100100100;
  urom[ 287] = 10'b0000000000;
  urom[ 288] = 10'b0000010111;
  urom[ 289] = 10'b0100101000;
  urom[ 290] = 10'b0000000000;
  urom[ 291] = 10'b0000010111;
  urom[ 292] = 10'b0100101100;
  urom[ 293] = 10'b0000000000;
  urom[ 294] = 10'b0000010111;
  urom[ 295] = 10'b0100110000;
  urom[ 296] = 10'b0011101110;
  urom[ 297] = 10'b0001100100;
  urom[ 298] = 10'b0100110100;
  urom[ 299] = 10'b0100111000;
  urom[ 300] = 10'b0100111100;
  urom[ 301] = 10'b0101000000;
  urom[ 302] = 10'b0101000100;
  urom[ 303] = 10'b0101001000;
  urom[ 304] = 10'b0101001100;
  urom[ 305] = 10'b0000010111;
  urom[ 306] = 10'b0000000100;
  urom[ 307] = 10'b0101010000;
  urom[ 308] = 10'b0101010100;
  urom[ 309] = 10'b0100111100;
  urom[ 310] = 10'b0101011000;
  urom[ 311] = 10'b0101001100;
  urom[ 312] = 10'b0000000000;
  urom[ 313] = 10'b0000000000;
  urom[ 314] = 10'b0000010111;
  urom[ 315] = 10'b0000000100;
  urom[ 316] = 10'b0101010000;
  urom[ 317] = 10'b0101010100;
  urom[ 318] = 10'b0100111100;
  urom[ 319] = 10'b0101011100;
  urom[ 320] = 10'b0101001100;
  urom[ 321] = 10'b0000000000;
  urom[ 322] = 10'b0000000000;
  urom[ 323] = 10'b0000010111;
  urom[ 324] = 10'b0000000100;
  urom[ 325] = 10'b0000001000;
  urom[ 326] = 10'b0000100000;
  urom[ 327] = 10'b0101100000;
  urom[ 328] = 10'b0101100100;
  urom[ 329] = 10'b0101101011;
  urom[ 330] = 10'b0101101110;
  urom[ 331] = 10'b0000000100;
  urom[ 332] = 10'b0000001000;
  urom[ 333] = 10'b0000100000;
  urom[ 334] = 10'b0000000100;
  urom[ 335] = 10'b0000001000;
  urom[ 336] = 10'b0101110000;
  urom[ 337] = 10'b0101110100;
  urom[ 338] = 10'b0000001100;
  urom[ 339] = 10'b0100100000;
  urom[ 340] = 10'b0101111000;
  urom[ 341] = 10'b0101111100;
  urom[ 342] = 10'b0110000011;
  urom[ 343] = 10'b0000000000;
  urom[ 344] = 10'b0000000000;
  urom[ 345] = 10'b0100100000;
  urom[ 346] = 10'b0101110100;
  urom[ 347] = 10'b0110000100;
  urom[ 348] = 10'b0100100000;
  urom[ 349] = 10'b0101111000;
  urom[ 350] = 10'b0110001000;
  urom[ 351] = 10'b0000010111;
  urom[ 352] = 10'b0110001100;
  urom[ 353] = 10'b0000001000;
  urom[ 354] = 10'b0110010000;
  urom[ 355] = 10'b0101110100;
  urom[ 356] = 10'b0000001100;
  urom[ 357] = 10'b0100100000;
  urom[ 358] = 10'b0101111000;
  urom[ 359] = 10'b0000001100;
  urom[ 360] = 10'b0110010100;
  urom[ 361] = 10'b0101100000;
  urom[ 362] = 10'b0110011000;
  urom[ 363] = 10'b0110011111;
  urom[ 364] = 10'b0000000000;
  urom[ 365] = 10'b0000000000;
  urom[ 366] = 10'b0100100000;
  urom[ 367] = 10'b0101110100;
  urom[ 368] = 10'b0000001100;
  urom[ 369] = 10'b0100100000;
  urom[ 370] = 10'b0101111000;
  urom[ 371] = 10'b0000001100;
  urom[ 372] = 10'b0110100000;
  urom[ 373] = 10'b0110100100;
  urom[ 374] = 10'b0110101000;
  urom[ 375] = 10'b0110101100;
  urom[ 376] = 10'b0110100100;
  urom[ 377] = 10'b0000001000;
  urom[ 378] = 10'b0101101011;
  urom[ 379] = 10'b0000000000;
  urom[ 380] = 10'b0000000000;
  urom[ 381] = 10'b0100100000;
  urom[ 382] = 10'b0110110000;
  urom[ 383] = 10'b0000001100;
  urom[ 384] = 10'b0100100000;
  urom[ 385] = 10'b0101110100;
  urom[ 386] = 10'b0000001100;
  urom[ 387] = 10'b0100100000;
  urom[ 388] = 10'b0101111000;
  urom[ 389] = 10'b0000001100;
  urom[ 390] = 10'b0110100000;
  urom[ 391] = 10'b0110110100;
  urom[ 392] = 10'b0000000000;
  urom[ 393] = 10'b0000000000;
  urom[ 394] = 10'b0110111000;
  urom[ 395] = 10'b0110111100;
  urom[ 396] = 10'b0000010111;
  urom[ 397] = 10'b0111000000;
  urom[ 398] = 10'b0111000100;
  urom[ 399] = 10'b0110101100;
  urom[ 400] = 10'b0111000000;
  urom[ 401] = 10'b0111000100;
  urom[ 402] = 10'b0101101011;
  urom[ 403] = 10'b0111000000;
  urom[ 404] = 10'b0111000100;
  urom[ 405] = 10'b0110101100;
  urom[ 406] = 10'b0111000000;
  urom[ 407] = 10'b0111000100;
  urom[ 408] = 10'b0111001011;
  urom[ 409] = 10'b0111000000;
  urom[ 410] = 10'b0111000100;
  urom[ 411] = 10'b0110101100;
  urom[ 412] = 10'b0111000000;
  urom[ 413] = 10'b0111000100;
  urom[ 414] = 10'b0111001100;
  urom[ 415] = 10'b0111000000;
  urom[ 416] = 10'b0111000100;
  urom[ 417] = 10'b0111010011;
  urom[ 418] = 10'b0000000100;
  urom[ 419] = 10'b0000001000;
  urom[ 420] = 10'b0000100000;
  urom[ 421] = 10'b0000100100;
  urom[ 422] = 10'b0111010100;
  urom[ 423] = 10'b0111011001;
  urom[ 424] = 10'b0111011110;
  urom[ 425] = 10'b0000010110;
  urom[ 426] = 10'b0000010110;
  urom[ 427] = 10'b0111100000;
  urom[ 428] = 10'b0111100100;
  urom[ 429] = 10'b0111101010;
  urom[ 430] = 10'b0111100000;
  urom[ 431] = 10'b0111101100;
  urom[ 432] = 10'b0111101010;
  urom[ 433] = 10'b0111110000;
  urom[ 434] = 10'b0111100100;
  urom[ 435] = 10'b0111110110;
  urom[ 436] = 10'b0111110000;
  urom[ 437] = 10'b0111101100;
  urom[ 438] = 10'b0111110110;
  urom[ 439] = 10'b0111100000;
  urom[ 440] = 10'b0111111000;
  urom[ 441] = 10'b0111101010;
  urom[ 442] = 10'b0111100000;
  urom[ 443] = 10'b0111111100;
  urom[ 444] = 10'b0111101010;
  urom[ 445] = 10'b0111110000;
  urom[ 446] = 10'b0111111000;
  urom[ 447] = 10'b0111110110;
  urom[ 448] = 10'b0111110000;
  urom[ 449] = 10'b0111111100;
  urom[ 450] = 10'b0111110110;
  urom[ 451] = 10'b0000000000;
  urom[ 452] = 10'b0000000000;
  urom[ 453] = 10'b0100100000;
  urom[ 454] = 10'b1000000000;
  urom[ 455] = 10'b0000001100;
  urom[ 456] = 10'b0100100000;
  urom[ 457] = 10'b1000000100;
  urom[ 458] = 10'b0000001100;
  urom[ 459] = 10'b0000010111;
  urom[ 460] = 10'b1000001000;
  urom[ 461] = 10'b0000001000;
  urom[ 462] = 10'b1000001100;
  urom[ 463] = 10'b1000001000;
  urom[ 464] = 10'b0000001000;
  urom[ 465] = 10'b1000010011;
  urom[ 466] = 10'b0000000000;
  urom[ 467] = 10'b0000000000;
  urom[ 468] = 10'b0100100000;
  urom[ 469] = 10'b1000010100;
  urom[ 470] = 10'b0000001100;
  urom[ 471] = 10'b0100100000;
  urom[ 472] = 10'b1000011000;
  urom[ 473] = 10'b0000001100;
  urom[ 474] = 10'b0000010111;
  urom[ 475] = 10'b1000001000;
  urom[ 476] = 10'b0000001000;
  urom[ 477] = 10'b0000110100;
  urom[ 478] = 10'b1000001000;
  urom[ 479] = 10'b0000001000;
  urom[ 480] = 10'b0000111011;
  urom[ 481] = 10'b0000000000;
  urom[ 482] = 10'b0000000000;
  urom[ 483] = 10'b0100100000;
  urom[ 484] = 10'b1000011100;
  urom[ 485] = 10'b0000001100;
  urom[ 486] = 10'b0100100000;
  urom[ 487] = 10'b1000100000;
  urom[ 488] = 10'b0000001100;
  urom[ 489] = 10'b0000010111;
  urom[ 490] = 10'b1000001000;
  urom[ 491] = 10'b0000001000;
  urom[ 492] = 10'b0000111100;
  urom[ 493] = 10'b1000001000;
  urom[ 494] = 10'b0000001000;
  urom[ 495] = 10'b0001000011;
  urom[ 496] = 10'b0000000000;
  urom[ 497] = 10'b0000000000;
  urom[ 498] = 10'b0100100000;
  urom[ 499] = 10'b1000100100;
  urom[ 500] = 10'b0000001100;
  urom[ 501] = 10'b0100100000;
  urom[ 502] = 10'b1000101000;
  urom[ 503] = 10'b0000001100;
  urom[ 504] = 10'b0000010111;
  urom[ 505] = 10'b1000001000;
  urom[ 506] = 10'b0000001000;
  urom[ 507] = 10'b0001000100;
  urom[ 508] = 10'b1000001000;
  urom[ 509] = 10'b0000001000;
  urom[ 510] = 10'b0001001011;
  urom[ 511] = 10'b1000101110;
  urom[ 512] = 10'b1000110010;
  urom[ 513] = 10'b1000110110;
  urom[ 514] = 10'b1000111010;
  urom[ 515] = 10'b1000111110;
  urom[ 516] = 10'b1001000010;
  urom[ 517] = 10'b1001000110;
  urom[ 518] = 10'b1001001010;
  urom[ 519] = 10'b1001001110;
  urom[ 520] = 10'b1001010010;
  urom[ 521] = 10'b0010000000;
  urom[ 522] = 10'b0000001000;
  urom[ 523] = 10'b0000100000;
  urom[ 524] = 10'b1001010100;
  urom[ 525] = 10'b0001101100;
  urom[ 526] = 10'b1001011000;
  urom[ 527] = 10'b1001011100;
  urom[ 528] = 10'b1001100000;
  urom[ 529] = 10'b1001100101;
  urom[ 530] = 10'b1001101010;
  urom[ 531] = 10'b0010000000;
  urom[ 532] = 10'b0000001000;
  urom[ 533] = 10'b0000100000;
  urom[ 534] = 10'b1001101100;
  urom[ 535] = 10'b1001011000;
  urom[ 536] = 10'b1001110000;
  urom[ 537] = 10'b1001011100;
  urom[ 538] = 10'b1001100000;
  urom[ 539] = 10'b1001100101;
  urom[ 540] = 10'b1001101010;
  urom[ 541] = 10'b1001110100;
  urom[ 542] = 10'b0000000000;
  urom[ 543] = 10'b0000010110;
  urom[ 544] = 10'b1001111000;
  urom[ 545] = 10'b0000000000;
  urom[ 546] = 10'b0000010110;
  urom[ 547] = 10'b1001111100;
  urom[ 548] = 10'b1010000000;
  urom[ 549] = 10'b1010000110;
  urom[ 550] = 10'b1001111100;
  urom[ 551] = 10'b1010001000;
  urom[ 552] = 10'b1010000110;
  urom[ 553] = 10'b1001111100;
  urom[ 554] = 10'b1010000000;
  urom[ 555] = 10'b1010001110;
  urom[ 556] = 10'b1001111100;
  urom[ 557] = 10'b1010010000;
  urom[ 558] = 10'b1010001110;
  urom[ 559] = 10'b1001111100;
  urom[ 560] = 10'b1010001000;
  urom[ 561] = 10'b1010001110;
  urom[ 562] = 10'b1001111100;
  urom[ 563] = 10'b1010010100;
  urom[ 564] = 10'b1010001110;
  urom[ 565] = 10'b0111100000;
  urom[ 566] = 10'b1010011000;
  urom[ 567] = 10'b0011100110;
  urom[ 568] = 10'b0111100000;
  urom[ 569] = 10'b1010011100;
  urom[ 570] = 10'b0011100110;
  urom[ 571] = 10'b0111100000;
  urom[ 572] = 10'b1010011000;
  urom[ 573] = 10'b0011101110;
  urom[ 574] = 10'b0111100000;
  urom[ 575] = 10'b1010100000;
  urom[ 576] = 10'b0011101110;
  urom[ 577] = 10'b0111100000;
  urom[ 578] = 10'b1010011100;
  urom[ 579] = 10'b0011101110;
  urom[ 580] = 10'b0111100000;
  urom[ 581] = 10'b1010100100;
  urom[ 582] = 10'b0011101110;
  urom[ 583] = 10'b1001111100;
  urom[ 584] = 10'b1010101000;
  urom[ 585] = 10'b1010101110;
  urom[ 586] = 10'b1001111100;
  urom[ 587] = 10'b1010110000;
  urom[ 588] = 10'b1010101110;
  urom[ 589] = 10'b1001111100;
  urom[ 590] = 10'b1010110100;
  urom[ 591] = 10'b1010101110;
  urom[ 592] = 10'b0111100000;
  urom[ 593] = 10'b1010111000;
  urom[ 594] = 10'b0010111010;
  urom[ 595] = 10'b0111100000;
  urom[ 596] = 10'b1010111100;
  urom[ 597] = 10'b0010111010;
  urom[ 598] = 10'b0111100000;
  urom[ 599] = 10'b1011000000;
  urom[ 600] = 10'b0010111010;
  urom[ 601] = 10'b1001111100;
  urom[ 602] = 10'b1011000100;
  urom[ 603] = 10'b0011000110;
  urom[ 604] = 10'b1001111100;
  urom[ 605] = 10'b1011001000;
  urom[ 606] = 10'b0011001110;
  urom[ 607] = 10'b1001111100;
  urom[ 608] = 10'b1011001000;
  urom[ 609] = 10'b0011011010;
  urom[ 610] = 10'b1001111100;
  urom[ 611] = 10'b1011001000;
  urom[ 612] = 10'b0011011110;
  urom[ 613] = 10'b0111100000;
  urom[ 614] = 10'b1011001100;
  urom[ 615] = 10'b0011000110;
  urom[ 616] = 10'b0111100000;
  urom[ 617] = 10'b1011010000;
  urom[ 618] = 10'b0011001110;
  urom[ 619] = 10'b0111100000;
  urom[ 620] = 10'b1010111000;
  urom[ 621] = 10'b0011010010;
  urom[ 622] = 10'b0111100000;
  urom[ 623] = 10'b1010111000;
  urom[ 624] = 10'b0011010110;
  urom[ 625] = 10'b0111100000;
  urom[ 626] = 10'b1011010000;
  urom[ 627] = 10'b0011011010;
  urom[ 628] = 10'b0111100000;
  urom[ 629] = 10'b1011010000;
  urom[ 630] = 10'b0011011110;
  urom[ 631] = 10'b1011010100;
  urom[ 632] = 10'b0000001000;
  urom[ 633] = 10'b0011100001;
  urom[ 634] = 10'b1010000110;
  urom[ 635] = 10'b1011010100;
  urom[ 636] = 10'b0000001000;
  urom[ 637] = 10'b0011101001;
  urom[ 638] = 10'b1010000110;
  urom[ 639] = 10'b1011010100;
  urom[ 640] = 10'b0000001000;
  urom[ 641] = 10'b0011100001;
  urom[ 642] = 10'b1010001110;
  urom[ 643] = 10'b1011010100;
  urom[ 644] = 10'b0000001000;
  urom[ 645] = 10'b0011110001;
  urom[ 646] = 10'b1010001110;
  urom[ 647] = 10'b1011010100;
  urom[ 648] = 10'b0000001000;
  urom[ 649] = 10'b0011101001;
  urom[ 650] = 10'b1010001110;
  urom[ 651] = 10'b1011010100;
  urom[ 652] = 10'b0000001000;
  urom[ 653] = 10'b0011110101;
  urom[ 654] = 10'b1010001110;
  urom[ 655] = 10'b1011010100;
  urom[ 656] = 10'b0000001000;
  urom[ 657] = 10'b0010101001;
  urom[ 658] = 10'b1010101110;
  urom[ 659] = 10'b1011010100;
  urom[ 660] = 10'b0000001000;
  urom[ 661] = 10'b0010111101;
  urom[ 662] = 10'b1010101110;
  urom[ 663] = 10'b1011010100;
  urom[ 664] = 10'b0000001000;
  urom[ 665] = 10'b0010110001;
  urom[ 666] = 10'b1010101110;
  urom[ 667] = 10'b1011011000;
  urom[ 668] = 10'b0000001000;
  urom[ 669] = 10'b0011100001;
  urom[ 670] = 10'b1011011110;
  urom[ 671] = 10'b1011011000;
  urom[ 672] = 10'b0000001000;
  urom[ 673] = 10'b0011101001;
  urom[ 674] = 10'b1011011110;
  urom[ 675] = 10'b1011011000;
  urom[ 676] = 10'b0000001000;
  urom[ 677] = 10'b0011100001;
  urom[ 678] = 10'b1011100010;
  urom[ 679] = 10'b1011011000;
  urom[ 680] = 10'b0000001000;
  urom[ 681] = 10'b0011110001;
  urom[ 682] = 10'b1011100010;
  urom[ 683] = 10'b1011011000;
  urom[ 684] = 10'b0000001000;
  urom[ 685] = 10'b0011101001;
  urom[ 686] = 10'b1011100010;
  urom[ 687] = 10'b1011011000;
  urom[ 688] = 10'b0000001000;
  urom[ 689] = 10'b0011110101;
  urom[ 690] = 10'b1011100010;
  urom[ 691] = 10'b1011011000;
  urom[ 692] = 10'b0000001000;
  urom[ 693] = 10'b0010101001;
  urom[ 694] = 10'b1011100110;
  urom[ 695] = 10'b1011011000;
  urom[ 696] = 10'b0000001000;
  urom[ 697] = 10'b0010111101;
  urom[ 698] = 10'b1011100110;
  urom[ 699] = 10'b1011011000;
  urom[ 700] = 10'b0000001000;
  urom[ 701] = 10'b0010110001;
  urom[ 702] = 10'b1011100110;
  urom[ 703] = 10'b1011010100;
  urom[ 704] = 10'b0000001000;
  urom[ 705] = 10'b0011000001;
  urom[ 706] = 10'b0011000110;
  urom[ 707] = 10'b1011010100;
  urom[ 708] = 10'b0000001000;
  urom[ 709] = 10'b0011001001;
  urom[ 710] = 10'b0011001110;
  urom[ 711] = 10'b1011010100;
  urom[ 712] = 10'b0000001000;
  urom[ 713] = 10'b0010101001;
  urom[ 714] = 10'b0011010010;
  urom[ 715] = 10'b1011010100;
  urom[ 716] = 10'b0000001000;
  urom[ 717] = 10'b0010101001;
  urom[ 718] = 10'b0011010110;
  urom[ 719] = 10'b1011010100;
  urom[ 720] = 10'b0000001000;
  urom[ 721] = 10'b0011001001;
  urom[ 722] = 10'b0011011010;
  urom[ 723] = 10'b1011010100;
  urom[ 724] = 10'b0000001000;
  urom[ 725] = 10'b0011001001;
  urom[ 726] = 10'b0011011110;
  urom[ 727] = 10'b1011011000;
  urom[ 728] = 10'b0000001000;
  urom[ 729] = 10'b0011000001;
  urom[ 730] = 10'b0011000110;
  urom[ 731] = 10'b1011011000;
  urom[ 732] = 10'b0000001000;
  urom[ 733] = 10'b0011001001;
  urom[ 734] = 10'b0011001110;
  urom[ 735] = 10'b1011011000;
  urom[ 736] = 10'b0000001000;
  urom[ 737] = 10'b0010101001;
  urom[ 738] = 10'b0011010010;
  urom[ 739] = 10'b1011011000;
  urom[ 740] = 10'b0000001000;
  urom[ 741] = 10'b0010101001;
  urom[ 742] = 10'b0011010110;
  urom[ 743] = 10'b1011011000;
  urom[ 744] = 10'b0000001000;
  urom[ 745] = 10'b0011001001;
  urom[ 746] = 10'b0011011010;
  urom[ 747] = 10'b1011011000;
  urom[ 748] = 10'b0000001000;
  urom[ 749] = 10'b0011001001;
  urom[ 750] = 10'b0011011110;
  urom[ 751] = 10'b0000000100;
  urom[ 752] = 10'b0000001000;
  urom[ 753] = 10'b0000100000;
  urom[ 754] = 10'b0000000100;
  urom[ 755] = 10'b0000001000;
  urom[ 756] = 10'b0001011100;
  urom[ 757] = 10'b0001110100;
  urom[ 758] = 10'b0000001000;
  urom[ 759] = 10'b0000011111;
  urom[ 760] = 10'b0000000100;
  urom[ 761] = 10'b0000001000;
  urom[ 762] = 10'b0000100000;
  urom[ 763] = 10'b0000000100;
  urom[ 764] = 10'b0000001000;
  urom[ 765] = 10'b0001011100;
  urom[ 766] = 10'b0001110100;
  urom[ 767] = 10'b0000001000;
  urom[ 768] = 10'b1011101000;
  urom[ 769] = 10'b0001111100;
  urom[ 770] = 10'b0000001000;
  urom[ 771] = 10'b0000110011;
  urom[ 772] = 10'b0000000100;
  urom[ 773] = 10'b0000001000;
  urom[ 774] = 10'b0000100000;
  urom[ 775] = 10'b0000000100;
  urom[ 776] = 10'b0000001000;
  urom[ 777] = 10'b0001011100;
  urom[ 778] = 10'b0001110100;
  urom[ 779] = 10'b0000001000;
  urom[ 780] = 10'b0001111000;
  urom[ 781] = 10'b0001111100;
  urom[ 782] = 10'b0000001000;
  urom[ 783] = 10'b0000111011;
  urom[ 784] = 10'b0000000100;
  urom[ 785] = 10'b0000001000;
  urom[ 786] = 10'b0000100000;
  urom[ 787] = 10'b0000000100;
  urom[ 788] = 10'b0000001000;
  urom[ 789] = 10'b0001011100;
  urom[ 790] = 10'b0001110100;
  urom[ 791] = 10'b0000001000;
  urom[ 792] = 10'b1011101100;
  urom[ 793] = 10'b0001111100;
  urom[ 794] = 10'b0000001000;
  urom[ 795] = 10'b0001000011;
  urom[ 796] = 10'b0000000100;
  urom[ 797] = 10'b0000001000;
  urom[ 798] = 10'b0000100000;
  urom[ 799] = 10'b0000000100;
  urom[ 800] = 10'b0000001000;
  urom[ 801] = 10'b0001011100;
  urom[ 802] = 10'b0001110100;
  urom[ 803] = 10'b0000001000;
  urom[ 804] = 10'b1011110000;
  urom[ 805] = 10'b0001111100;
  urom[ 806] = 10'b0000001000;
  urom[ 807] = 10'b0001001011;
  urom[ 808] = 10'b0000000100;
  urom[ 809] = 10'b1011110100;
  urom[ 810] = 10'b0000100000;
  urom[ 811] = 10'b0000000100;
  urom[ 812] = 10'b0000001000;
  urom[ 813] = 10'b0001011100;
  urom[ 814] = 10'b0001110100;
  urom[ 815] = 10'b0000001100;
  urom[ 816] = 10'b0000010111;
  urom[ 817] = 10'b0000000100;
  urom[ 818] = 10'b0000001000;
  urom[ 819] = 10'b0000100000;
  urom[ 820] = 10'b0000000100;
  urom[ 821] = 10'b1011111000;
  urom[ 822] = 10'b0001011100;
  urom[ 823] = 10'b0001110100;
  urom[ 824] = 10'b0000001100;
  urom[ 825] = 10'b1011111100;
  urom[ 826] = 10'b1100000000;
  urom[ 827] = 10'b0000001100;
  urom[ 828] = 10'b0000010111;
  urom[ 829] = 10'b0000000100;
  urom[ 830] = 10'b0000001000;
  urom[ 831] = 10'b0000100000;
  urom[ 832] = 10'b0000000100;
  urom[ 833] = 10'b1100000100;
  urom[ 834] = 10'b0001011100;
  urom[ 835] = 10'b0001110100;
  urom[ 836] = 10'b0000001100;
  urom[ 837] = 10'b1011111100;
  urom[ 838] = 10'b1100001000;
  urom[ 839] = 10'b0000001100;
  urom[ 840] = 10'b0000010111;
  urom[ 841] = 10'b0000000100;
  urom[ 842] = 10'b0000001000;
  urom[ 843] = 10'b0000100000;
  urom[ 844] = 10'b0000000100;
  urom[ 845] = 10'b1100001100;
  urom[ 846] = 10'b0001011100;
  urom[ 847] = 10'b0001110100;
  urom[ 848] = 10'b0000001100;
  urom[ 849] = 10'b1011111100;
  urom[ 850] = 10'b1100010000;
  urom[ 851] = 10'b0000001100;
  urom[ 852] = 10'b0000010111;
  urom[ 853] = 10'b0000000100;
  urom[ 854] = 10'b0000001000;
  urom[ 855] = 10'b0000100000;
  urom[ 856] = 10'b0000000100;
  urom[ 857] = 10'b1100010100;
  urom[ 858] = 10'b0001011100;
  urom[ 859] = 10'b0001110100;
  urom[ 860] = 10'b0000001100;
  urom[ 861] = 10'b1011111100;
  urom[ 862] = 10'b1100011000;
  urom[ 863] = 10'b0000001100;
  urom[ 864] = 10'b0000010111;
  urom[ 865] = 10'b0001001100;
  urom[ 866] = 10'b1100011100;
  urom[ 867] = 10'b0011100001;
  urom[ 868] = 10'b0011100110;
  urom[ 869] = 10'b0001001100;
  urom[ 870] = 10'b1100011100;
  urom[ 871] = 10'b0011101001;
  urom[ 872] = 10'b0011100110;
  urom[ 873] = 10'b0001001100;
  urom[ 874] = 10'b1100011100;
  urom[ 875] = 10'b0011100001;
  urom[ 876] = 10'b0011101110;
  urom[ 877] = 10'b0001001100;
  urom[ 878] = 10'b1100011100;
  urom[ 879] = 10'b0011110001;
  urom[ 880] = 10'b0011101110;
  urom[ 881] = 10'b0001001100;
  urom[ 882] = 10'b1100011100;
  urom[ 883] = 10'b0011101001;
  urom[ 884] = 10'b0011101110;
  urom[ 885] = 10'b0001001100;
  urom[ 886] = 10'b1100011100;
  urom[ 887] = 10'b0011110101;
  urom[ 888] = 10'b0011101110;
  urom[ 889] = 10'b0001001100;
  urom[ 890] = 10'b1100011100;
  urom[ 891] = 10'b0010101001;
  urom[ 892] = 10'b0010111010;
  urom[ 893] = 10'b0001001100;
  urom[ 894] = 10'b1100011100;
  urom[ 895] = 10'b0010111101;
  urom[ 896] = 10'b0010111010;
  urom[ 897] = 10'b0001001100;
  urom[ 898] = 10'b1100011100;
  urom[ 899] = 10'b0010110001;
  urom[ 900] = 10'b0010111010;
  urom[ 901] = 10'b0001001100;
  urom[ 902] = 10'b1100011100;
  urom[ 903] = 10'b0011000001;
  urom[ 904] = 10'b0011000110;
  urom[ 905] = 10'b0001001100;
  urom[ 906] = 10'b1100011100;
  urom[ 907] = 10'b0011001001;
  urom[ 908] = 10'b0011001110;
  urom[ 909] = 10'b0001001100;
  urom[ 910] = 10'b1100011100;
  urom[ 911] = 10'b0010101001;
  urom[ 912] = 10'b0011010010;
  urom[ 913] = 10'b0001001100;
  urom[ 914] = 10'b1100011100;
  urom[ 915] = 10'b0010101001;
  urom[ 916] = 10'b0011010110;
  urom[ 917] = 10'b0001001100;
  urom[ 918] = 10'b1100011100;
  urom[ 919] = 10'b0011001001;
  urom[ 920] = 10'b0011011010;
  urom[ 921] = 10'b0001001100;
  urom[ 922] = 10'b1100011100;
  urom[ 923] = 10'b0011001001;
  urom[ 924] = 10'b0011011110;
  urom[ 925] = 10'b0000000100;
  urom[ 926] = 10'b0000001000;
  urom[ 927] = 10'b0000100000;
  urom[ 928] = 10'b1100100000;
  urom[ 929] = 10'b0000001000;
  urom[ 930] = 10'b0011100001;
  urom[ 931] = 10'b0011100110;
  urom[ 932] = 10'b0000000100;
  urom[ 933] = 10'b0000001000;
  urom[ 934] = 10'b0000100000;
  urom[ 935] = 10'b1100100000;
  urom[ 936] = 10'b0000001000;
  urom[ 937] = 10'b0011101001;
  urom[ 938] = 10'b0011100110;
  urom[ 939] = 10'b0000000100;
  urom[ 940] = 10'b0000001000;
  urom[ 941] = 10'b0000100000;
  urom[ 942] = 10'b1100100000;
  urom[ 943] = 10'b0000001000;
  urom[ 944] = 10'b0011100001;
  urom[ 945] = 10'b0011101110;
  urom[ 946] = 10'b0000000100;
  urom[ 947] = 10'b0000001000;
  urom[ 948] = 10'b0000100000;
  urom[ 949] = 10'b1100100000;
  urom[ 950] = 10'b0000001000;
  urom[ 951] = 10'b0011110001;
  urom[ 952] = 10'b0011101110;
  urom[ 953] = 10'b0000000100;
  urom[ 954] = 10'b0000001000;
  urom[ 955] = 10'b0000100000;
  urom[ 956] = 10'b1100100000;
  urom[ 957] = 10'b0000001000;
  urom[ 958] = 10'b0011101001;
  urom[ 959] = 10'b0011101110;
  urom[ 960] = 10'b0000000100;
  urom[ 961] = 10'b0000001000;
  urom[ 962] = 10'b0000100000;
  urom[ 963] = 10'b1100100000;
  urom[ 964] = 10'b0000001000;
  urom[ 965] = 10'b0011110101;
  urom[ 966] = 10'b0011101110;
  urom[ 967] = 10'b0000000100;
  urom[ 968] = 10'b0000001000;
  urom[ 969] = 10'b0000100000;
  urom[ 970] = 10'b1100100000;
  urom[ 971] = 10'b0000001000;
  urom[ 972] = 10'b0010101001;
  urom[ 973] = 10'b0010111010;
  urom[ 974] = 10'b0000000100;
  urom[ 975] = 10'b0000001000;
  urom[ 976] = 10'b0000100000;
  urom[ 977] = 10'b1100100000;
  urom[ 978] = 10'b0000001000;
  urom[ 979] = 10'b0010111101;
  urom[ 980] = 10'b0010111010;
  urom[ 981] = 10'b0000000100;
  urom[ 982] = 10'b0000001000;
  urom[ 983] = 10'b0000100000;
  urom[ 984] = 10'b1100100000;
  urom[ 985] = 10'b0000001000;
  urom[ 986] = 10'b0010110001;
  urom[ 987] = 10'b0010111010;
  urom[ 988] = 10'b0000000100;
  urom[ 989] = 10'b0000001000;
  urom[ 990] = 10'b0000100000;
  urom[ 991] = 10'b1100100000;
  urom[ 992] = 10'b0000001000;
  urom[ 993] = 10'b0011000001;
  urom[ 994] = 10'b0011000110;
  urom[ 995] = 10'b0000000100;
  urom[ 996] = 10'b0000001000;
  urom[ 997] = 10'b0000100000;
  urom[ 998] = 10'b1100100000;
  urom[ 999] = 10'b0000001000;
  urom[1000] = 10'b0011001001;
  urom[1001] = 10'b0011001110;
  urom[1002] = 10'b0000000100;
  urom[1003] = 10'b0000001000;
  urom[1004] = 10'b0000100000;
  urom[1005] = 10'b1100100000;
  urom[1006] = 10'b0000001000;
  urom[1007] = 10'b0010101001;
  urom[1008] = 10'b0011010010;
  urom[1009] = 10'b0000000100;
  urom[1010] = 10'b0000001000;
  urom[1011] = 10'b0000100000;
  urom[1012] = 10'b1100100000;
  urom[1013] = 10'b0000001000;
  urom[1014] = 10'b0010101001;
  urom[1015] = 10'b0011010110;
  urom[1016] = 10'b0000000100;
  urom[1017] = 10'b0000001000;
  urom[1018] = 10'b0000100000;
  urom[1019] = 10'b1100100000;
  urom[1020] = 10'b0000001000;
  urom[1021] = 10'b0011001001;
  urom[1022] = 10'b0011011010;
  urom[1023] = 10'b0000000100;
  urom[1024] = 10'b0000001000;
  urom[1025] = 10'b0000100000;
  urom[1026] = 10'b1100100000;
  urom[1027] = 10'b0000001000;
  urom[1028] = 10'b0011001001;
  urom[1029] = 10'b0011011110;
end
