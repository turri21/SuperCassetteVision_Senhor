s_nc nrom [201];
initial begin
  nrom[   0] = 54'b000000000000000000000000000000000000000000000000000000;
  nrom[   1] = 54'b000000000000000000000000001001000000000000000000000000;
  nrom[   2] = 54'b000000000000000000000000000000100000000000000000000000;
  nrom[   3] = 54'b000000000000000000000000000000010000000000000000000000;
  nrom[   4] = 54'b000110100010010001000000000000000000000000000000000000;
  nrom[   5] = 54'b000000000000000000000000000000000000000000000000000001;
  nrom[   6] = 54'b000000111010010001000000000000000000000000000000000000;
  nrom[   7] = 54'b000000011010100001000000000000000000000000000000000001;
  nrom[   8] = 54'b000000011100100001000000000000000000000000000000000000;
  nrom[   9] = 54'b000000000000000000010100000001000000000000000000000000;
  nrom[  10] = 54'b000000000010100001000000000000000000000000000000000001;
  nrom[  11] = 54'b000000010010100001000000000000000000000000000000000000;
  nrom[  12] = 54'b000000010100100001000000000000000000000000000000000001;
  nrom[  13] = 54'b000000000110100001000000000000000000000000000000000000;
  nrom[  14] = 54'b000000000100100001000000000000000000000000000000000001;
  nrom[  15] = 54'b000000001010100001000000000000000000000000000000000000;
  nrom[  16] = 54'b000000001000100001000000000000000000000000000000000001;
  nrom[  17] = 54'b000000001110100001000000000000000000000000000000000000;
  nrom[  18] = 54'b000000001100100001000000000000000000000000000000000001;
  nrom[  19] = 54'b000000000000000000011101110001000000000000000000000010;
  nrom[  20] = 54'b000000100000010010011101110001000000000000000000000010;
  nrom[  21] = 54'b000111000000010010011101110001000000000000000000000010;
  nrom[  22] = 54'b000000100000010010010100000001000000000000000000000000;
  nrom[  23] = 54'b000000000000100011000000000000000001001000000000000000;
  nrom[  24] = 54'b000000000000110010010100000001000000000000000000000000;
  nrom[  25] = 54'b000101100000010011000000000000000000000000000000000000;
  nrom[  26] = 54'b000000100000010100000000000000000001010000000000000000;
  nrom[  27] = 54'b000000011100110001000000000000000000000000000000000000;
  nrom[  28] = 54'b000110000000010011000000000000000001101000000000000000;
  nrom[  29] = 54'b000000000000110000011000000001000000000000000000000000;
  nrom[  30] = 54'b000000000110100001100000000000000000000000000000000000;
  nrom[  31] = 54'b000000000000000000100100000101000000000000000000000000;
  nrom[  32] = 54'b000000000000000000010000000001000000000000000000000000;
  nrom[  33] = 54'b000000000000000000010001000100100000000000000000000000;
  nrom[  34] = 54'b000111000000010010001100000001000000000000000000000000;
  nrom[  35] = 54'b000000000000000000001100110100010000000000000000000000;
  nrom[  36] = 54'b000001100000010011000000000000000100000000000000000000;
  nrom[  37] = 54'b000000000110110001000000000000000000000000000000000000;
  nrom[  38] = 54'b000000000000000000000000000010000000000000000100000001;
  nrom[  39] = 54'b000000000000001000000000000000000000000000000000000001;
  nrom[  40] = 54'b000000000100001000000000000000000000000000000000000001;
  nrom[  41] = 54'b000000000000100011000000000000000000000000000000000000;
  nrom[  42] = 54'b000000000000100100000000000000000110000000000000000000;
  nrom[  43] = 54'b000000000000000000000000000000000000000010000000000001;
  nrom[  44] = 54'b000000000000100100000000000000000101000000000000000000;
  nrom[  45] = 54'b000000100000010011000000001001000000000000000000000000;
  nrom[  46] = 54'b000000000010110001000000000000000000000010000000000001;
  nrom[  47] = 54'b000000000000100100000000000000000111000000000000000000;
  nrom[  48] = 54'b000000000000100100000000000000000010010100000000000000;
  nrom[  49] = 54'b000000000000000000000000000000000000000011100110000001;
  nrom[  50] = 54'b000000000000100100000000000000000010000100000000000000;
  nrom[  51] = 54'b000000000000000000000000000000000000000011100100000001;
  nrom[  52] = 54'b000000000000000000000000000000000000000010001010000001;
  nrom[  53] = 54'b000000000000000000000000000000000000000010001000000001;
  nrom[  54] = 54'b000000000000000000000000000000000000000011101010000001;
  nrom[  55] = 54'b000000000000000000000000000000000000000011101000000001;
  nrom[  56] = 54'b000000000000100100000000000000000001000000000000000000;
  nrom[  57] = 54'b000000000010110001000000000000000000000011100110000001;
  nrom[  58] = 54'b000000000000100100000000000000000010000100000000000000;
  nrom[  59] = 54'b000000000010110001000000000000000000000011100000000001;
  nrom[  60] = 54'b000000000000100100000000000000000001110000000000000000;
  nrom[  61] = 54'b000000000000100100000000000000000010110100000000000000;
  nrom[  62] = 54'b000000000000100011000000000000000011000000000000000000;
  nrom[  63] = 54'b000000000000000000000000000000000000000010100100000001;
  nrom[  64] = 54'b000000000000100011000000000000000100000000000000000000;
  nrom[  65] = 54'b000110100000010011000000000000000011000000000000000000;
  nrom[  66] = 54'b000000011010110001000000000000000000000010100100000001;
  nrom[  67] = 54'b000110100000010011000000000000000100000000000000000000;
  nrom[  68] = 54'b000000000000000000000100010100000000000000000000000000;
  nrom[  69] = 54'b000000000000000000001000100100000000000000000000000000;
  nrom[  70] = 54'b000000000000000000001100110100000000000000000000000000;
  nrom[  71] = 54'b000000000000000000010001000100000000000000000000000000;
  nrom[  72] = 54'b000000000000000000000100010010000000000000000000000000;
  nrom[  73] = 54'b000000000000000000001000100010000000000000000000000000;
  nrom[  74] = 54'b000000000000000000001100110010000000000000000000000000;
  nrom[  75] = 54'b000000000000000000010001000010000000000000000000000000;
  nrom[  76] = 54'b000000100000010011000000000000000001000000000000000100;
  nrom[  77] = 54'b000000000001010100000000000000000000000000000000000000;
  nrom[  78] = 54'b000000000000000000000000000000000001000000000000000000;
  nrom[  79] = 54'b000000010110110001000000000000000000000000000000000000;
  nrom[  80] = 54'b000110000000010011000000000000000000000000000000000000;
  nrom[  81] = 54'b000000000001010100000000000000000000000000000000001000;
  nrom[  82] = 54'b000000000000000000000000000000000001100000000000000000;
  nrom[  83] = 54'b000000011000110001000000000000000000000000000000000000;
  nrom[  84] = 54'b000101100000010011000000000000100000000000000000000000;
  nrom[  85] = 54'b000000000000100100000000000000000001000000000000000000;
  nrom[  86] = 54'b000110000000010011000000000000000001101000000000000000;
  nrom[  87] = 54'b000110000000010011000000000000000001101100000000000000;
  nrom[  88] = 54'b000000000000000000000000000001000000000000000000000000;
  nrom[  89] = 54'b000111010110010001000000000000100000000000000000000000;
  nrom[  90] = 54'b000000011000100001000000000000000000000000000000000001;
  nrom[  91] = 54'b000000000000000000001000000111000000000000000000000001;
  nrom[  92] = 54'b000000000000100011000100010010000001001000000000000000;
  nrom[  93] = 54'b000110000000010010000100000001000000000000000000000000;
  nrom[  94] = 54'b000101100000010010000100000001000000000000000000000000;
  nrom[  95] = 54'b000111010110010001000000000000010000000000000000000000;
  nrom[  96] = 54'b000000011000110001000000000000000000000000000000000001;
  nrom[  97] = 54'b000001011000010001000000000000010000000000000000000000;
  nrom[  98] = 54'b000001110110010001000000000000010000000000000000000000;
  nrom[  99] = 54'b000000000000000000000000001000000000000000000000000000;
  nrom[ 100] = 54'b000000011100100001000100010010000000000000000000000000;
  nrom[ 101] = 54'b000000000000000000000000000010000000000000000000000000;
  nrom[ 102] = 54'b000000011001010001000000000000100000000000000000010000;
  nrom[ 103] = 54'b000000010110100001000000000000000000000000000000000001;
  nrom[ 104] = 54'b000000011101010001000000000000000000000000000000011000;
  nrom[ 105] = 54'b000000000000000000011000000001000000000000000000000000;
  nrom[ 106] = 54'b001000011101010001000000000000100000000000000000011000;
  nrom[ 107] = 54'b000000010110100001000000000000000000000000000000000000;
  nrom[ 108] = 54'b000100000000010010000100000001000000000000000000000000;
  nrom[ 109] = 54'b000000011000000001000000000000000000000000000000000000;
  nrom[ 110] = 54'b000000010111010001000000000000000000000000000000100000;
  nrom[ 111] = 54'b000000000000000000000000000000000000000000010000000000;
  nrom[ 112] = 54'b000000000000000000000100000001000000000000000000000000;
  nrom[ 113] = 54'b000000000000000000000100010100100000000000000000000000;
  nrom[ 114] = 54'b000000011000100001000000000000000000000000000010000001;
  nrom[ 115] = 54'b000000011000100001000000000000000000000000000000000000;
  nrom[ 116] = 54'b000000010000100001000000000000000000000000000000000001;
  nrom[ 117] = 54'b000000000001010100000000000000100000000000000000101000;
  nrom[ 118] = 54'b000000000000100011000000000000000110000000000000000000;
  nrom[ 119] = 54'b000000000000000000000000000000000000000000001010000001;
  nrom[ 120] = 54'b000000100000010011000000000000000000000000000000000000;
  nrom[ 121] = 54'b000000000000000000000000000000001001110000000000000000;
  nrom[ 122] = 54'b000000000010110001000000000000000000000001000000000001;
  nrom[ 123] = 54'b000000000000000000000000000000001011110000000000000000;
  nrom[ 124] = 54'b000001100000010011000000000000000000000000000000000000;
  nrom[ 125] = 54'b000000000110110001000000000000000000000001000000000001;
  nrom[ 126] = 54'b000000000000000000000000000000001000000000000000000000;
  nrom[ 127] = 54'b000000000000000000000000000000001010000000000000000000;
  nrom[ 128] = 54'b000000000000010010000100000001000000000000000000000000;
  nrom[ 129] = 54'b000000100000010010000100000001000000000000000000000000;
  nrom[ 130] = 54'b000000000000000000000100010101000000000000000000000000;
  nrom[ 131] = 54'b000000000010100001000000000000000000000000000000000000;
  nrom[ 132] = 54'b000000000000100001000000000000000000000000000000000001;
  nrom[ 133] = 54'b000001000000010010000100000001000000000000000000000000;
  nrom[ 134] = 54'b000001100000010010000100000001000000000000000000000000;
  nrom[ 135] = 54'b000010000000010010000100000001000000000000000000000000;
  nrom[ 136] = 54'b000010100000010010000100000001000000000000000000000000;
  nrom[ 137] = 54'b000011000000010010000100000001000000000000000000000000;
  nrom[ 138] = 54'b000011100000010010000100000001000000000000000000000000;
  nrom[ 139] = 54'b000000000000000000000000000000000000000000001100000001;
  nrom[ 140] = 54'b000000000000000000000000000000000000000000010010000001;
  nrom[ 141] = 54'b000000000000000000000000000000000000000000010110000001;
  nrom[ 142] = 54'b000000000000000000000000000000000000000000001110000001;
  nrom[ 143] = 54'b000000000000000000000000000000000000000000010100000001;
  nrom[ 144] = 54'b000000000000000000000000000000000000000000011000000001;
  nrom[ 145] = 54'b001000000000000101000000000000000000000000000000000001;
  nrom[ 146] = 54'b000000000000000101000000000000000000000000000000000001;
  nrom[ 147] = 54'b000000000000000111000000000000000000000000000000000001;
  nrom[ 148] = 54'b001000000000000111000000000000000000000000000000000001;
  nrom[ 149] = 54'b000111000000010011000000000000001110000000000000000000;
  nrom[ 150] = 54'b000000100000010011000000000000001100000000000000000000;
  nrom[ 151] = 54'b000111000000110010010000000001000000000000000000000000;
  nrom[ 152] = 54'b000111000000010011000000000000011100000000000000000000;
  nrom[ 153] = 54'b000000100000010011000000000000001101000000000000000000;
  nrom[ 154] = 54'b000000000010110001000000000000000000000000000000000001;
  nrom[ 155] = 54'b000111000000010011000000000000001101000000000000000000;
  nrom[ 156] = 54'b000000000000110011000000000000001110000000000000000000;
  nrom[ 157] = 54'b000000000011000001000000000000000000000000000001000000;
  nrom[ 158] = 54'b000000100000010110000000000000000000000000000001000000;
  nrom[ 159] = 54'b000110100000010011000000000000000000000000000000000000;
  nrom[ 160] = 54'b000000100000010100000000000000000001000000000000000000;
  nrom[ 161] = 54'b000000011010110001000000000000000000000011100110000001;
  nrom[ 162] = 54'b000000100000010100000000000000000010000100000000000000;
  nrom[ 163] = 54'b000000011010110001000000000000000000000011100000000001;
  nrom[ 164] = 54'b000000100000010100000000000000000001110000000000000000;
  nrom[ 165] = 54'b000000100000010100000000000000000010110100000000000000;
  nrom[ 166] = 54'b000110100000010100000000000000000001000000000000000000;
  nrom[ 167] = 54'b000110100000010100000000000000000010000100000000000000;
  nrom[ 168] = 54'b000110100000010100000000000000000001110000000000000000;
  nrom[ 169] = 54'b000110100000010100000000000000000010110100000000000000;
  nrom[ 170] = 54'b000000100000010100000000000000000110000000000000000000;
  nrom[ 171] = 54'b000000011010110001000000000000000000000010000000000001;
  nrom[ 172] = 54'b000000100000010100000000000000000111000000000000000000;
  nrom[ 173] = 54'b000000100000010100000000000000000101000000000000000000;
  nrom[ 174] = 54'b000110100000010100000000000000000110000000000000000000;
  nrom[ 175] = 54'b000110100000010100000000000000000111000000000000000000;
  nrom[ 176] = 54'b000110100000010100000000000000000101000000000000000000;
  nrom[ 177] = 54'b000000100000010100000000000000000010010100000000000000;
  nrom[ 178] = 54'b000000100000010100000000000000000010000100000000000000;
  nrom[ 179] = 54'b000110100000010100000000000000000010010100000000000000;
  nrom[ 180] = 54'b000110100000010100000000000000000010000100000000000000;
  nrom[ 181] = 54'b000110100000010011000000001001000000000000000000000000;
  nrom[ 182] = 54'b000000000001000011000000001001000000000000000000000000;
  nrom[ 183] = 54'b000000000000110110000000000000000000000011100110000001;
  nrom[ 184] = 54'b000000000000110110000000000000000000000011100000000001;
  nrom[ 185] = 54'b000000000000110110000000000000000000000010000000000001;
  nrom[ 186] = 54'b000000010010100001100000000000000000000000000000000000;
  nrom[ 187] = 54'b000000001010100001100000000000000000000000000000000000;
  nrom[ 188] = 54'b000000001110100001100000000000000000000000000000000000;
  nrom[ 189] = 54'b000110100000010010000000000000100000000000000000000000;
  nrom[ 190] = 54'b000100100000010010000000000000100000000000000000000000;
  nrom[ 191] = 54'b000000000000000000100000000000000000000000000000000000;
  nrom[ 192] = 54'b000101000000010010100100000101000000000000000000000000;
  nrom[ 193] = 54'b000001100000010010000000000000100000000000000000000000;
  nrom[ 194] = 54'b000001000000010010100100000101000000000000000000000000;
  nrom[ 195] = 54'b000010100000010010000000000000100000000000000000000000;
  nrom[ 196] = 54'b000010000000010010100100000101000000000000000000000000;
  nrom[ 197] = 54'b000011100000010010000000000000100000000000000000000000;
  nrom[ 198] = 54'b000011000000010010100100000101000000000000000000000000;
  nrom[ 199] = 54'b000000100000010011000000000000100000000000000000000000;
  nrom[ 200] = 54'b000000100000010011010100000001000000000000000000000000;
end
