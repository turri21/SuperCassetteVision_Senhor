// NEC uPD7800 testbench: reset
//
// Copyright (c) 2024 David Hunter
//
// This program is GPL licensed. See COPYING for the full license.

`timescale 1us / 1ns

module reset_tb();

reg         clk, res;
reg         cp1p, cp1n, cp2p, cp2n;
reg [7:0]   din;

wire [15:0] a;
wire [7:0]  dout;

initial begin
  $timeformat(-6, 0, " us", 1);

  $dumpfile("tb/reset_tb.vcd");
  $dumpvars();
end

upd7800 dut
  (
   .CLK(clk),
   .CP1_POSEDGE(cp1p),
   .CP1_NEGEDGE(cp1n),
   .CP2_POSEDGE(cp2p),
   .CP2_NEGEDGE(cp2n),
   .RESETB(~res),
   .A(a),
   .DB_I(8'hzz),
   .DB_O(),
   .DB_OE(),
   .M1()
   );


initial begin
  cp1p = 0;
  cp1n = 0;
  cp2p = 0;
  cp2n = 0;
  res = 1;
  clk = 1;
end

initial forever begin :ckgen
  #0.125 clk = ~clk;
end

initial forever begin :cpgen
  @(posedge clk) cp2n <= 0; cp1p <= 1;
  @(posedge clk) cp1p <= 0; cp1n <= 1;
  @(posedge clk) cp1n <= 0; cp2p <= 1;
  @(posedge clk) cp2p <= 0; cp2n <= 1;
end

wire cp2 = dut.cp2;

initial #0 begin
  #11 @(posedge clk) ;
  res = 0;
  #11 @(posedge clk) ;

  $finish;
end


endmodule

// Local Variables:
// compile-command: "cd .. && iverilog -g2012 -grelative-include -s reset_tb -o reset_tb.vvp upd7800.sv tb/reset_tb.sv && tb/reset_tb.vvp"
// End:
