s_uc urom [582];
initial begin
  urom[   0] = 11'b00000000010;
  urom[   1] = 11'b00000001000;
  urom[   2] = 11'b00000010000;
  urom[   3] = 11'b00000000000;
  urom[   4] = 11'b00000001000;
  urom[   5] = 11'b00000010000;
  urom[   6] = 11'b00000000011;
  urom[   7] = 11'b00000100000;
  urom[   8] = 11'b00000000000;
  urom[   9] = 11'b00000000010;
  urom[  10] = 11'b00000101000;
  urom[  11] = 11'b00000000000;
  urom[  12] = 11'b00000000010;
  urom[  13] = 11'b00000001000;
  urom[  14] = 11'b00000010000;
  urom[  15] = 11'b00000110011;
  urom[  16] = 11'b00000001000;
  urom[  17] = 11'b00000010000;
  urom[  18] = 11'b00000111000;
  urom[  19] = 11'b00001000000;
  urom[  20] = 11'b00000010000;
  urom[  21] = 11'b00001001011;
  urom[  22] = 11'b00000001000;
  urom[  23] = 11'b00000010000;
  urom[  24] = 11'b00001010000;
  urom[  25] = 11'b00000001000;
  urom[  26] = 11'b00000010000;
  urom[  27] = 11'b00001011011;
  urom[  28] = 11'b00000001000;
  urom[  29] = 11'b00000010000;
  urom[  30] = 11'b00001100000;
  urom[  31] = 11'b00000001000;
  urom[  32] = 11'b00000010000;
  urom[  33] = 11'b00001101011;
  urom[  34] = 11'b00000001000;
  urom[  35] = 11'b00000010000;
  urom[  36] = 11'b00001110000;
  urom[  37] = 11'b00000001000;
  urom[  38] = 11'b00000010000;
  urom[  39] = 11'b00001111011;
  urom[  40] = 11'b00000001000;
  urom[  41] = 11'b00000010000;
  urom[  42] = 11'b00010000000;
  urom[  43] = 11'b00000001000;
  urom[  44] = 11'b00000010000;
  urom[  45] = 11'b00010001011;
  urom[  46] = 11'b00010010000;
  urom[  47] = 11'b00000010000;
  urom[  48] = 11'b00001001011;
  urom[  49] = 11'b00010011000;
  urom[  50] = 11'b00000011000;
  urom[  51] = 11'b00000000011;
  urom[  52] = 11'b00000001000;
  urom[  53] = 11'b00000010000;
  urom[  54] = 11'b00000111000;
  urom[  55] = 11'b00010100000;
  urom[  56] = 11'b00000011000;
  urom[  57] = 11'b00000000011;
  urom[  58] = 11'b00000001000;
  urom[  59] = 11'b00000010000;
  urom[  60] = 11'b00000111000;
  urom[  61] = 11'b00010101000;
  urom[  62] = 11'b00000011000;
  urom[  63] = 11'b00000000011;
  urom[  64] = 11'b00000001000;
  urom[  65] = 11'b00000010000;
  urom[  66] = 11'b00000111000;
  urom[  67] = 11'b00000001000;
  urom[  68] = 11'b00000010000;
  urom[  69] = 11'b00010110000;
  urom[  70] = 11'b00010111000;
  urom[  71] = 11'b00000011000;
  urom[  72] = 11'b00000000011;
  urom[  73] = 11'b00011000000;
  urom[  74] = 11'b00000000000;
  urom[  75] = 11'b00000000000;
  urom[  76] = 11'b00011001000;
  urom[  77] = 11'b00011010000;
  urom[  78] = 11'b00000000000;
  urom[  79] = 11'b00011011000;
  urom[  80] = 11'b00000000000;
  urom[  81] = 11'b00000000000;
  urom[  82] = 11'b00011100000;
  urom[  83] = 11'b00000010000;
  urom[  84] = 11'b00011101000;
  urom[  85] = 11'b00011110000;
  urom[  86] = 11'b00000010000;
  urom[  87] = 11'b00001101011;
  urom[  88] = 11'b00011111000;
  urom[  89] = 11'b00100000000;
  urom[  90] = 11'b00000111000;
  urom[  91] = 11'b00100001000;
  urom[  92] = 11'b00100010000;
  urom[  93] = 11'b00000000000;
  urom[  94] = 11'b00100011000;
  urom[  95] = 11'b00100100000;
  urom[  96] = 11'b00100101011;
  urom[  97] = 11'b00000001000;
  urom[  98] = 11'b00000010000;
  urom[  99] = 11'b00000111000;
  urom[ 100] = 11'b00001000000;
  urom[ 101] = 11'b00000010000;
  urom[ 102] = 11'b00100110000;
  urom[ 103] = 11'b00000001000;
  urom[ 104] = 11'b00000010000;
  urom[ 105] = 11'b00100111000;
  urom[ 106] = 11'b00010111000;
  urom[ 107] = 11'b00000011000;
  urom[ 108] = 11'b00101000011;
  urom[ 109] = 11'b00000001000;
  urom[ 110] = 11'b00000010000;
  urom[ 111] = 11'b00000111000;
  urom[ 112] = 11'b00001000000;
  urom[ 113] = 11'b00000010000;
  urom[ 114] = 11'b00100110000;
  urom[ 115] = 11'b00000001000;
  urom[ 116] = 11'b00000010000;
  urom[ 117] = 11'b00101001000;
  urom[ 118] = 11'b00010111000;
  urom[ 119] = 11'b00000011000;
  urom[ 120] = 11'b00101000011;
  urom[ 121] = 11'b00101010000;
  urom[ 122] = 11'b00000010000;
  urom[ 123] = 11'b00100111001;
  urom[ 124] = 11'b00101011010;
  urom[ 125] = 11'b00101010000;
  urom[ 126] = 11'b00000010000;
  urom[ 127] = 11'b00101100001;
  urom[ 128] = 11'b00101011010;
  urom[ 129] = 11'b00101010000;
  urom[ 130] = 11'b00000010000;
  urom[ 131] = 11'b00101001001;
  urom[ 132] = 11'b00101011010;
  urom[ 133] = 11'b00000001000;
  urom[ 134] = 11'b00000010000;
  urom[ 135] = 11'b00000111000;
  urom[ 136] = 11'b00001000000;
  urom[ 137] = 11'b00000010000;
  urom[ 138] = 11'b00100110000;
  urom[ 139] = 11'b00000001000;
  urom[ 140] = 11'b00000010000;
  urom[ 141] = 11'b00100111001;
  urom[ 142] = 11'b00101101010;
  urom[ 143] = 11'b00000001000;
  urom[ 144] = 11'b00000010000;
  urom[ 145] = 11'b00000111000;
  urom[ 146] = 11'b00001000000;
  urom[ 147] = 11'b00000010000;
  urom[ 148] = 11'b00100110000;
  urom[ 149] = 11'b00000001000;
  urom[ 150] = 11'b00000010000;
  urom[ 151] = 11'b00101110001;
  urom[ 152] = 11'b00101111010;
  urom[ 153] = 11'b00000001000;
  urom[ 154] = 11'b00110000000;
  urom[ 155] = 11'b00101110001;
  urom[ 156] = 11'b00110001010;
  urom[ 157] = 11'b00000001000;
  urom[ 158] = 11'b00110000000;
  urom[ 159] = 11'b00101110001;
  urom[ 160] = 11'b00110010010;
  urom[ 161] = 11'b00000001000;
  urom[ 162] = 11'b00110000000;
  urom[ 163] = 11'b00100111001;
  urom[ 164] = 11'b00101101010;
  urom[ 165] = 11'b00000001000;
  urom[ 166] = 11'b00110000000;
  urom[ 167] = 11'b00100111001;
  urom[ 168] = 11'b00110011010;
  urom[ 169] = 11'b00000001000;
  urom[ 170] = 11'b00110000000;
  urom[ 171] = 11'b00101110001;
  urom[ 172] = 11'b00101111010;
  urom[ 173] = 11'b00000001000;
  urom[ 174] = 11'b00110000000;
  urom[ 175] = 11'b00101110001;
  urom[ 176] = 11'b00110100010;
  urom[ 177] = 11'b00101010000;
  urom[ 178] = 11'b00000010000;
  urom[ 179] = 11'b00110101001;
  urom[ 180] = 11'b00110110010;
  urom[ 181] = 11'b00101010000;
  urom[ 182] = 11'b00000010000;
  urom[ 183] = 11'b00101110001;
  urom[ 184] = 11'b00110111010;
  urom[ 185] = 11'b00101010000;
  urom[ 186] = 11'b00000010000;
  urom[ 187] = 11'b00110101001;
  urom[ 188] = 11'b00111000010;
  urom[ 189] = 11'b00101010000;
  urom[ 190] = 11'b00000010000;
  urom[ 191] = 11'b00111001001;
  urom[ 192] = 11'b00111000010;
  urom[ 193] = 11'b00101010000;
  urom[ 194] = 11'b00000010000;
  urom[ 195] = 11'b00101110001;
  urom[ 196] = 11'b00111000010;
  urom[ 197] = 11'b00101010000;
  urom[ 198] = 11'b00000010000;
  urom[ 199] = 11'b00111010001;
  urom[ 200] = 11'b00111000010;
  urom[ 201] = 11'b00000001000;
  urom[ 202] = 11'b00000010000;
  urom[ 203] = 11'b00000111000;
  urom[ 204] = 11'b00001000000;
  urom[ 205] = 11'b00000010000;
  urom[ 206] = 11'b00111011000;
  urom[ 207] = 11'b00010111000;
  urom[ 208] = 11'b00000011000;
  urom[ 209] = 11'b00110001011;
  urom[ 210] = 11'b00000001000;
  urom[ 211] = 11'b00000010000;
  urom[ 212] = 11'b00000111000;
  urom[ 213] = 11'b00001000000;
  urom[ 214] = 11'b00000010000;
  urom[ 215] = 11'b00111100000;
  urom[ 216] = 11'b00010111000;
  urom[ 217] = 11'b00000011000;
  urom[ 218] = 11'b00110010011;
  urom[ 219] = 11'b00111101000;
  urom[ 220] = 11'b00111110010;
  urom[ 221] = 11'b00111111000;
  urom[ 222] = 11'b01000000010;
  urom[ 223] = 11'b01000001000;
  urom[ 224] = 11'b00000000000;
  urom[ 225] = 11'b00000000011;
  urom[ 226] = 11'b01000010000;
  urom[ 227] = 11'b00000000000;
  urom[ 228] = 11'b00000000011;
  urom[ 229] = 11'b01000011000;
  urom[ 230] = 11'b00000000000;
  urom[ 231] = 11'b00000000011;
  urom[ 232] = 11'b01000100000;
  urom[ 233] = 11'b00000000000;
  urom[ 234] = 11'b00000000011;
  urom[ 235] = 11'b01000101000;
  urom[ 236] = 11'b00000000000;
  urom[ 237] = 11'b00000000011;
  urom[ 238] = 11'b01000110000;
  urom[ 239] = 11'b00000000000;
  urom[ 240] = 11'b00000000011;
  urom[ 241] = 11'b01000111000;
  urom[ 242] = 11'b00000000000;
  urom[ 243] = 11'b00000000011;
  urom[ 244] = 11'b01001000000;
  urom[ 245] = 11'b00000000000;
  urom[ 246] = 11'b00000000011;
  urom[ 247] = 11'b01001001000;
  urom[ 248] = 11'b00111000010;
  urom[ 249] = 11'b00011000000;
  urom[ 250] = 11'b01001010000;
  urom[ 251] = 11'b01001011000;
  urom[ 252] = 11'b01001100000;
  urom[ 253] = 11'b01001101000;
  urom[ 254] = 11'b01001110000;
  urom[ 255] = 11'b01001111000;
  urom[ 256] = 11'b01010000000;
  urom[ 257] = 11'b00000000011;
  urom[ 258] = 11'b00000001000;
  urom[ 259] = 11'b01010001000;
  urom[ 260] = 11'b01010010000;
  urom[ 261] = 11'b01001100000;
  urom[ 262] = 11'b01010011000;
  urom[ 263] = 11'b01010000000;
  urom[ 264] = 11'b00000000000;
  urom[ 265] = 11'b00000000000;
  urom[ 266] = 11'b00000000011;
  urom[ 267] = 11'b00000001000;
  urom[ 268] = 11'b01010001000;
  urom[ 269] = 11'b01010010000;
  urom[ 270] = 11'b01001100000;
  urom[ 271] = 11'b01010100000;
  urom[ 272] = 11'b01010000000;
  urom[ 273] = 11'b00000000000;
  urom[ 274] = 11'b00000000000;
  urom[ 275] = 11'b00000000011;
  urom[ 276] = 11'b00000001000;
  urom[ 277] = 11'b00000010000;
  urom[ 278] = 11'b00000111000;
  urom[ 279] = 11'b01010101000;
  urom[ 280] = 11'b01010110000;
  urom[ 281] = 11'b01010111011;
  urom[ 282] = 11'b01011000010;
  urom[ 283] = 11'b01011001000;
  urom[ 284] = 11'b00000010000;
  urom[ 285] = 11'b01011010000;
  urom[ 286] = 11'b01011011000;
  urom[ 287] = 11'b00000011000;
  urom[ 288] = 11'b01000101000;
  urom[ 289] = 11'b01011100000;
  urom[ 290] = 11'b00000011000;
  urom[ 291] = 11'b01011101000;
  urom[ 292] = 11'b01010101000;
  urom[ 293] = 11'b01011110000;
  urom[ 294] = 11'b01011111011;
  urom[ 295] = 11'b00000000000;
  urom[ 296] = 11'b00000000000;
  urom[ 297] = 11'b01000101000;
  urom[ 298] = 11'b01011011000;
  urom[ 299] = 11'b00000011000;
  urom[ 300] = 11'b01000101000;
  urom[ 301] = 11'b01011100000;
  urom[ 302] = 11'b00000011000;
  urom[ 303] = 11'b01100000000;
  urom[ 304] = 11'b01100001000;
  urom[ 305] = 11'b01100010000;
  urom[ 306] = 11'b01011111000;
  urom[ 307] = 11'b01100001000;
  urom[ 308] = 11'b00000010000;
  urom[ 309] = 11'b01010111011;
  urom[ 310] = 11'b00000000000;
  urom[ 311] = 11'b00000000000;
  urom[ 312] = 11'b01000101000;
  urom[ 313] = 11'b01100011000;
  urom[ 314] = 11'b00000011000;
  urom[ 315] = 11'b01000101000;
  urom[ 316] = 11'b01011011000;
  urom[ 317] = 11'b00000011000;
  urom[ 318] = 11'b01000101000;
  urom[ 319] = 11'b01011100000;
  urom[ 320] = 11'b00000011000;
  urom[ 321] = 11'b01100000000;
  urom[ 322] = 11'b01100100000;
  urom[ 323] = 11'b00000000000;
  urom[ 324] = 11'b00000000000;
  urom[ 325] = 11'b01100101000;
  urom[ 326] = 11'b01100110000;
  urom[ 327] = 11'b00000000011;
  urom[ 328] = 11'b01100111000;
  urom[ 329] = 11'b01101000000;
  urom[ 330] = 11'b01011111000;
  urom[ 331] = 11'b01100111000;
  urom[ 332] = 11'b01101000000;
  urom[ 333] = 11'b01010111011;
  urom[ 334] = 11'b01100111000;
  urom[ 335] = 11'b01101000000;
  urom[ 336] = 11'b01011111000;
  urom[ 337] = 11'b01100111000;
  urom[ 338] = 11'b01101000000;
  urom[ 339] = 11'b01010111000;
  urom[ 340] = 11'b01100111000;
  urom[ 341] = 11'b01101000000;
  urom[ 342] = 11'b01101001011;
  urom[ 343] = 11'b00000001000;
  urom[ 344] = 11'b00000010000;
  urom[ 345] = 11'b00000111000;
  urom[ 346] = 11'b00001000000;
  urom[ 347] = 11'b01101010000;
  urom[ 348] = 11'b01101011001;
  urom[ 349] = 11'b01101100010;
  urom[ 350] = 11'b00000000010;
  urom[ 351] = 11'b01101101000;
  urom[ 352] = 11'b01101110000;
  urom[ 353] = 11'b01101111010;
  urom[ 354] = 11'b01101101000;
  urom[ 355] = 11'b01110000000;
  urom[ 356] = 11'b01101111010;
  urom[ 357] = 11'b01110001000;
  urom[ 358] = 11'b01101110000;
  urom[ 359] = 11'b01110010010;
  urom[ 360] = 11'b01110001000;
  urom[ 361] = 11'b01110000000;
  urom[ 362] = 11'b01110010010;
  urom[ 363] = 11'b01101101000;
  urom[ 364] = 11'b01110011000;
  urom[ 365] = 11'b01101111010;
  urom[ 366] = 11'b01101101000;
  urom[ 367] = 11'b01110100000;
  urom[ 368] = 11'b01101111010;
  urom[ 369] = 11'b01110001000;
  urom[ 370] = 11'b01110011000;
  urom[ 371] = 11'b01110010010;
  urom[ 372] = 11'b01110001000;
  urom[ 373] = 11'b01110100000;
  urom[ 374] = 11'b01110010010;
  urom[ 375] = 11'b00000000000;
  urom[ 376] = 11'b00000000000;
  urom[ 377] = 11'b01000101000;
  urom[ 378] = 11'b01110101000;
  urom[ 379] = 11'b00000011000;
  urom[ 380] = 11'b01000101000;
  urom[ 381] = 11'b01110110000;
  urom[ 382] = 11'b00000011000;
  urom[ 383] = 11'b00000000011;
  urom[ 384] = 11'b01110111000;
  urom[ 385] = 11'b00000010000;
  urom[ 386] = 11'b00001001000;
  urom[ 387] = 11'b01110111000;
  urom[ 388] = 11'b00000010000;
  urom[ 389] = 11'b01111000011;
  urom[ 390] = 11'b00000000000;
  urom[ 391] = 11'b00000000000;
  urom[ 392] = 11'b01000101000;
  urom[ 393] = 11'b01111001000;
  urom[ 394] = 11'b00000011000;
  urom[ 395] = 11'b01000101000;
  urom[ 396] = 11'b01111010000;
  urom[ 397] = 11'b00000011000;
  urom[ 398] = 11'b00000000011;
  urom[ 399] = 11'b01110111000;
  urom[ 400] = 11'b00000010000;
  urom[ 401] = 11'b00001100000;
  urom[ 402] = 11'b01110111000;
  urom[ 403] = 11'b00000010000;
  urom[ 404] = 11'b00001101011;
  urom[ 405] = 11'b00000000000;
  urom[ 406] = 11'b00000000000;
  urom[ 407] = 11'b01000101000;
  urom[ 408] = 11'b01111011000;
  urom[ 409] = 11'b00000011000;
  urom[ 410] = 11'b01000101000;
  urom[ 411] = 11'b01111100000;
  urom[ 412] = 11'b00000011000;
  urom[ 413] = 11'b00000000011;
  urom[ 414] = 11'b01110111000;
  urom[ 415] = 11'b00000010000;
  urom[ 416] = 11'b00001110000;
  urom[ 417] = 11'b01110111000;
  urom[ 418] = 11'b00000010000;
  urom[ 419] = 11'b00001111011;
  urom[ 420] = 11'b00000000000;
  urom[ 421] = 11'b00000000000;
  urom[ 422] = 11'b01000101000;
  urom[ 423] = 11'b01111101000;
  urom[ 424] = 11'b00000011000;
  urom[ 425] = 11'b01000101000;
  urom[ 426] = 11'b01111110000;
  urom[ 427] = 11'b00000011000;
  urom[ 428] = 11'b00000000011;
  urom[ 429] = 11'b01110111000;
  urom[ 430] = 11'b00000010000;
  urom[ 431] = 11'b00010000000;
  urom[ 432] = 11'b01110111000;
  urom[ 433] = 11'b00000010000;
  urom[ 434] = 11'b00010001011;
  urom[ 435] = 11'b01111111010;
  urom[ 436] = 11'b10000000010;
  urom[ 437] = 11'b10000001010;
  urom[ 438] = 11'b10000010010;
  urom[ 439] = 11'b10000011010;
  urom[ 440] = 11'b10000100010;
  urom[ 441] = 11'b10000101000;
  urom[ 442] = 11'b00000000000;
  urom[ 443] = 11'b00000000010;
  urom[ 444] = 11'b10000110000;
  urom[ 445] = 11'b00000000000;
  urom[ 446] = 11'b00000000010;
  urom[ 447] = 11'b10000111000;
  urom[ 448] = 11'b10001000000;
  urom[ 449] = 11'b01000000010;
  urom[ 450] = 11'b10000111000;
  urom[ 451] = 11'b10001001000;
  urom[ 452] = 11'b00111110010;
  urom[ 453] = 11'b10000111000;
  urom[ 454] = 11'b10001000000;
  urom[ 455] = 11'b10001010010;
  urom[ 456] = 11'b10000111000;
  urom[ 457] = 11'b10001011000;
  urom[ 458] = 11'b10001010010;
  urom[ 459] = 11'b10000111000;
  urom[ 460] = 11'b10001001000;
  urom[ 461] = 11'b10001010010;
  urom[ 462] = 11'b10000111000;
  urom[ 463] = 11'b10001100000;
  urom[ 464] = 11'b10001010010;
  urom[ 465] = 11'b01101101000;
  urom[ 466] = 11'b10001101000;
  urom[ 467] = 11'b00110110010;
  urom[ 468] = 11'b01101101000;
  urom[ 469] = 11'b10001110000;
  urom[ 470] = 11'b00110111010;
  urom[ 471] = 11'b01101101000;
  urom[ 472] = 11'b10001101000;
  urom[ 473] = 11'b00111000010;
  urom[ 474] = 11'b01101101000;
  urom[ 475] = 11'b10001111000;
  urom[ 476] = 11'b00111000010;
  urom[ 477] = 11'b01101101000;
  urom[ 478] = 11'b10001110000;
  urom[ 479] = 11'b00111000010;
  urom[ 480] = 11'b01101101000;
  urom[ 481] = 11'b10010000000;
  urom[ 482] = 11'b00111000010;
  urom[ 483] = 11'b10010001000;
  urom[ 484] = 11'b00000010000;
  urom[ 485] = 11'b00110101001;
  urom[ 486] = 11'b01000000010;
  urom[ 487] = 11'b10010001000;
  urom[ 488] = 11'b00000010000;
  urom[ 489] = 11'b00101110001;
  urom[ 490] = 11'b00111110010;
  urom[ 491] = 11'b10010001000;
  urom[ 492] = 11'b00000010000;
  urom[ 493] = 11'b00110101001;
  urom[ 494] = 11'b10001010010;
  urom[ 495] = 11'b10010001000;
  urom[ 496] = 11'b00000010000;
  urom[ 497] = 11'b00111001001;
  urom[ 498] = 11'b10001010010;
  urom[ 499] = 11'b00000001000;
  urom[ 500] = 11'b10010010000;
  urom[ 501] = 11'b00100111001;
  urom[ 502] = 11'b00110011010;
  urom[ 503] = 11'b10010001000;
  urom[ 504] = 11'b00000010000;
  urom[ 505] = 11'b00101110001;
  urom[ 506] = 11'b10001010010;
  urom[ 507] = 11'b10010001000;
  urom[ 508] = 11'b00000010000;
  urom[ 509] = 11'b00111010001;
  urom[ 510] = 11'b10001010010;
  urom[ 511] = 11'b10010011000;
  urom[ 512] = 11'b00000010000;
  urom[ 513] = 11'b00100111001;
  urom[ 514] = 11'b10010100010;
  urom[ 515] = 11'b10010011000;
  urom[ 516] = 11'b00000010000;
  urom[ 517] = 11'b00101100001;
  urom[ 518] = 11'b10010100010;
  urom[ 519] = 11'b10010011000;
  urom[ 520] = 11'b00000010000;
  urom[ 521] = 11'b00101001001;
  urom[ 522] = 11'b10010100010;
  urom[ 523] = 11'b00000001000;
  urom[ 524] = 11'b10010010000;
  urom[ 525] = 11'b00100111001;
  urom[ 526] = 11'b00101101010;
  urom[ 527] = 11'b00000001000;
  urom[ 528] = 11'b10010101000;
  urom[ 529] = 11'b00100111001;
  urom[ 530] = 11'b00101101010;
  urom[ 531] = 11'b00000001000;
  urom[ 532] = 11'b10010101000;
  urom[ 533] = 11'b00100111001;
  urom[ 534] = 11'b00110011010;
  urom[ 535] = 11'b00000001000;
  urom[ 536] = 11'b00000010000;
  urom[ 537] = 11'b00000111000;
  urom[ 538] = 11'b00000001000;
  urom[ 539] = 11'b00000010000;
  urom[ 540] = 11'b00010110000;
  urom[ 541] = 11'b00011100000;
  urom[ 542] = 11'b00000010000;
  urom[ 543] = 11'b00000110011;
  urom[ 544] = 11'b00000001000;
  urom[ 545] = 11'b10010110000;
  urom[ 546] = 11'b00000111000;
  urom[ 547] = 11'b00000001000;
  urom[ 548] = 11'b00000010000;
  urom[ 549] = 11'b00010110000;
  urom[ 550] = 11'b00011100000;
  urom[ 551] = 11'b00000011000;
  urom[ 552] = 11'b00000000011;
  urom[ 553] = 11'b00010010000;
  urom[ 554] = 11'b00110000000;
  urom[ 555] = 11'b00110101001;
  urom[ 556] = 11'b00111000010;
  urom[ 557] = 11'b00010010000;
  urom[ 558] = 11'b00110000000;
  urom[ 559] = 11'b00101110001;
  urom[ 560] = 11'b00111000010;
  urom[ 561] = 11'b00000001000;
  urom[ 562] = 11'b00000010000;
  urom[ 563] = 11'b00000111000;
  urom[ 564] = 11'b10010111000;
  urom[ 565] = 11'b00000010000;
  urom[ 566] = 11'b00110101001;
  urom[ 567] = 11'b00111000010;
  urom[ 568] = 11'b00000001000;
  urom[ 569] = 11'b00000010000;
  urom[ 570] = 11'b00000111000;
  urom[ 571] = 11'b10010111000;
  urom[ 572] = 11'b00000010000;
  urom[ 573] = 11'b00100111001;
  urom[ 574] = 11'b00101011010;
  urom[ 575] = 11'b00000001000;
  urom[ 576] = 11'b00000010000;
  urom[ 577] = 11'b00000111000;
  urom[ 578] = 11'b10010111000;
  urom[ 579] = 11'b00000010000;
  urom[ 580] = 11'b00101001000;
  urom[ 581] = 11'b00101011010;
end
