    ird_lut['h00a] = {UA_MOV_A_RF_IR210, 1'd1, 2'd0};
    ird_lut['h00b] = {UA_MOV_A_RF_IR210, 1'd1, 2'd0};
    ird_lut['h00c] = {UA_MOV_A_RF_IR210, 1'd1, 2'd0};
    ird_lut['h00d] = {UA_MOV_A_RF_IR210, 1'd1, 2'd0};
    ird_lut['h00e] = {UA_MOV_A_RF_IR210, 1'd1, 2'd0};
    ird_lut['h00f] = {UA_MOV_A_RF_IR210, 1'd1, 2'd0};
    ird_lut['h01a] = {UA_MOV_RF_IR210_A, 1'd1, 2'd0};
    ird_lut['h01b] = {UA_MOV_RF_IR210_A, 1'd1, 2'd0};
    ird_lut['h01c] = {UA_MOV_RF_IR210_A, 1'd1, 2'd0};
    ird_lut['h01d] = {UA_MOV_RF_IR210_A, 1'd1, 2'd0};
    ird_lut['h01e] = {UA_MOV_RF_IR210_A, 1'd1, 2'd0};
    ird_lut['h01f] = {UA_MOV_RF_IR210_A, 1'd1, 2'd0};
    ird_lut['h068] = {UA_MOV_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h069] = {UA_MOV_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h06a] = {UA_MOV_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h06b] = {UA_MOV_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h06c] = {UA_MOV_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h06d] = {UA_MOV_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h06e] = {UA_MOV_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h06f] = {UA_MOV_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h028] = {UA_LD_A_WA, 1'd0, 2'd1};
    ird_lut['h004] = {UA_LDX_SP_IMM, 1'd0, 2'd2};
    ird_lut['h014] = {UA_LDX_BC_IMM, 1'd0, 2'd2};
    ird_lut['h024] = {UA_LDX_DE_IMM, 1'd0, 2'd2};
    ird_lut['h034] = {UA_LDX_HL_IMM, 1'd0, 2'd2};
    ird_lut['h029] = {UA_LDAX, 1'd0, 2'd0};
    ird_lut['h02a] = {UA_LDAX, 1'd0, 2'd0};
    ird_lut['h02b] = {UA_LDAX, 1'd0, 2'd0};
    ird_lut['h02c] = {UA_LDAX, 1'd0, 2'd0};
    ird_lut['h02d] = {UA_LDAX, 1'd0, 2'd0};
    ird_lut['h02e] = {UA_LDAX, 1'd0, 2'd0};
    ird_lut['h02f] = {UA_LDAX, 1'd0, 2'd0};
    ird_lut['h03a] = {UA_STX_A, 1'd0, 2'd0};
    ird_lut['h03b] = {UA_STX_A, 1'd0, 2'd0};
    ird_lut['h03c] = {UA_STX_A, 1'd0, 2'd0};
    ird_lut['h03d] = {UA_STX_A, 1'd0, 2'd0};
    ird_lut['h048] = {UA_STX_RF_W, 1'd0, 2'd1};
    ird_lut['h049] = {UA_STX_RF_W, 1'd0, 2'd1};
    ird_lut['h04a] = {UA_STX_RF_W, 1'd0, 2'd1};
    ird_lut['h04b] = {UA_STX_RF_W, 1'd0, 2'd1};
    ird_lut['h038] = {UA_STW_A, 1'd0, 2'd1};
    ird_lut['h071] = {UA_STW_IMM, 1'd0, 2'd2};
    ird_lut['h021] = {UA_TABLE, 1'd0, 2'd0};
    ird_lut['h031] = {UA_BLOCK, 1'd0, 2'd0};
    ird_lut['h005] = {UA_AND_WA_IMM, 1'd0, 2'd2};
    ird_lut['h015] = {UA_OR_WA_IMM, 1'd0, 2'd2};
    ird_lut['h007] = {UA_AND_A_IMM, 1'd0, 2'd1};
    ird_lut['h016] = {UA_XOR_A_IMM, 1'd0, 2'd1};
    ird_lut['h017] = {UA_OR_A_IMM, 1'd0, 2'd1};
    ird_lut['h045] = {UA_ON_WA_IMM, 1'd0, 2'd1};
    ird_lut['h065] = {UA_NEQ_WA_IMM, 1'd0, 2'd1};
    ird_lut['h027] = {UA_GT_A_IMM, 1'd0, 2'd1};
    ird_lut['h037] = {UA_LT_A_IMM, 1'd0, 2'd1};
    ird_lut['h047] = {UA_ON_A_IMM, 1'd0, 2'd1};
    ird_lut['h057] = {UA_OFF_A_IMM, 1'd0, 2'd1};
    ird_lut['h067] = {UA_NEQ_A_IMM, 1'd0, 2'd1};
    ird_lut['h077] = {UA_EQ_A_IMM, 1'd0, 2'd1};
    ird_lut['h026] = {UA_ADDNC_A_IMM, 1'd0, 2'd1};
    ird_lut['h036] = {UA_SUBNB_A_IMM, 1'd0, 2'd1};
    ird_lut['h046] = {UA_ADD_A_IMM, 1'd0, 2'd1};
    ird_lut['h056] = {UA_ADC_A_IMM, 1'd0, 2'd1};
    ird_lut['h066] = {UA_SUB_A_IMM, 1'd0, 2'd1};
    ird_lut['h076] = {UA_SBB_A_IMM, 1'd0, 2'd1};
    ird_lut['h020] = {UA_INCR_WA, 1'd0, 2'd0};
    ird_lut['h030] = {UA_DECR_WA, 1'd0, 2'd0};
    ird_lut['h041] = {UA_INCR_RF_IR210, 1'd1, 2'd0};
    ird_lut['h042] = {UA_INCR_RF_IR210, 1'd1, 2'd0};
    ird_lut['h043] = {UA_INCR_RF_IR210, 1'd1, 2'd0};
    ird_lut['h051] = {UA_DECR_RF_IR210, 1'd1, 2'd0};
    ird_lut['h052] = {UA_DECR_RF_IR210, 1'd1, 2'd0};
    ird_lut['h053] = {UA_DECR_RF_IR210, 1'd1, 2'd0};
    ird_lut['h002] = {UA_INC_SP, 1'd0, 2'd0};
    ird_lut['h012] = {UA_INC_BC, 1'd0, 2'd0};
    ird_lut['h022] = {UA_INC_DE, 1'd0, 2'd0};
    ird_lut['h032] = {UA_INC_HL, 1'd0, 2'd0};
    ird_lut['h003] = {UA_DEC_SP, 1'd0, 2'd0};
    ird_lut['h013] = {UA_DEC_BC, 1'd0, 2'd0};
    ird_lut['h023] = {UA_DEC_DE, 1'd0, 2'd0};
    ird_lut['h033] = {UA_DEC_HL, 1'd0, 2'd0};
    ird_lut['h061] = {UA_DAA, 1'd1, 2'd0};
    ird_lut['h0c0] = {UA_JR, 1'd0, 2'd0};
    ird_lut['h0c1] = {UA_JR, 1'd0, 2'd0};
    ird_lut['h0c2] = {UA_JR, 1'd0, 2'd0};
    ird_lut['h0c3] = {UA_JR, 1'd0, 2'd0};
    ird_lut['h0c4] = {UA_JR, 1'd0, 2'd0};
    ird_lut['h0c5] = {UA_JR, 1'd0, 2'd0};
    ird_lut['h0c6] = {UA_JR, 1'd0, 2'd0};
    ird_lut['h0c7] = {UA_JR, 1'd0, 2'd0};
    ird_lut['h0c8] = {UA_JR, 1'd0, 2'd0};
    ird_lut['h0c9] = {UA_JR, 1'd0, 2'd0};
    ird_lut['h0ca] = {UA_JR, 1'd0, 2'd0};
    ird_lut['h0cb] = {UA_JR, 1'd0, 2'd0};
    ird_lut['h0cc] = {UA_JR, 1'd0, 2'd0};
    ird_lut['h0cd] = {UA_JR, 1'd0, 2'd0};
    ird_lut['h0ce] = {UA_JR, 1'd0, 2'd0};
    ird_lut['h0cf] = {UA_JR, 1'd0, 2'd0};
    ird_lut['h0d0] = {UA_JR, 1'd0, 2'd0};
    ird_lut['h0d1] = {UA_JR, 1'd0, 2'd0};
    ird_lut['h0d2] = {UA_JR, 1'd0, 2'd0};
    ird_lut['h0d3] = {UA_JR, 1'd0, 2'd0};
    ird_lut['h0d4] = {UA_JR, 1'd0, 2'd0};
    ird_lut['h0d5] = {UA_JR, 1'd0, 2'd0};
    ird_lut['h0d6] = {UA_JR, 1'd0, 2'd0};
    ird_lut['h0d7] = {UA_JR, 1'd0, 2'd0};
    ird_lut['h0d8] = {UA_JR, 1'd0, 2'd0};
    ird_lut['h0d9] = {UA_JR, 1'd0, 2'd0};
    ird_lut['h0da] = {UA_JR, 1'd0, 2'd0};
    ird_lut['h0db] = {UA_JR, 1'd0, 2'd0};
    ird_lut['h0dc] = {UA_JR, 1'd0, 2'd0};
    ird_lut['h0dd] = {UA_JR, 1'd0, 2'd0};
    ird_lut['h0de] = {UA_JR, 1'd0, 2'd0};
    ird_lut['h0df] = {UA_JR, 1'd0, 2'd0};
    ird_lut['h0e0] = {UA_JR, 1'd0, 2'd0};
    ird_lut['h0e1] = {UA_JR, 1'd0, 2'd0};
    ird_lut['h0e2] = {UA_JR, 1'd0, 2'd0};
    ird_lut['h0e3] = {UA_JR, 1'd0, 2'd0};
    ird_lut['h0e4] = {UA_JR, 1'd0, 2'd0};
    ird_lut['h0e5] = {UA_JR, 1'd0, 2'd0};
    ird_lut['h0e6] = {UA_JR, 1'd0, 2'd0};
    ird_lut['h0e7] = {UA_JR, 1'd0, 2'd0};
    ird_lut['h0e8] = {UA_JR, 1'd0, 2'd0};
    ird_lut['h0e9] = {UA_JR, 1'd0, 2'd0};
    ird_lut['h0ea] = {UA_JR, 1'd0, 2'd0};
    ird_lut['h0eb] = {UA_JR, 1'd0, 2'd0};
    ird_lut['h0ec] = {UA_JR, 1'd0, 2'd0};
    ird_lut['h0ed] = {UA_JR, 1'd0, 2'd0};
    ird_lut['h0ee] = {UA_JR, 1'd0, 2'd0};
    ird_lut['h0ef] = {UA_JR, 1'd0, 2'd0};
    ird_lut['h0f0] = {UA_JR, 1'd0, 2'd0};
    ird_lut['h0f1] = {UA_JR, 1'd0, 2'd0};
    ird_lut['h0f2] = {UA_JR, 1'd0, 2'd0};
    ird_lut['h0f3] = {UA_JR, 1'd0, 2'd0};
    ird_lut['h0f4] = {UA_JR, 1'd0, 2'd0};
    ird_lut['h0f5] = {UA_JR, 1'd0, 2'd0};
    ird_lut['h0f6] = {UA_JR, 1'd0, 2'd0};
    ird_lut['h0f7] = {UA_JR, 1'd0, 2'd0};
    ird_lut['h0f8] = {UA_JR, 1'd0, 2'd0};
    ird_lut['h0f9] = {UA_JR, 1'd0, 2'd0};
    ird_lut['h0fa] = {UA_JR, 1'd0, 2'd0};
    ird_lut['h0fb] = {UA_JR, 1'd0, 2'd0};
    ird_lut['h0fc] = {UA_JR, 1'd0, 2'd0};
    ird_lut['h0fd] = {UA_JR, 1'd0, 2'd0};
    ird_lut['h0fe] = {UA_JR, 1'd0, 2'd0};
    ird_lut['h0ff] = {UA_JR, 1'd0, 2'd0};
    ird_lut['h04e] = {UA_JRE_P, 1'd0, 2'd1};
    ird_lut['h04f] = {UA_JRE_N, 1'd0, 2'd1};
    ird_lut['h054] = {UA_JMP, 1'd0, 2'd2};
    ird_lut['h073] = {UA_JB, 1'd1, 2'd0};
    ird_lut['h078] = {UA_CALF, 1'd0, 2'd1};
    ird_lut['h079] = {UA_CALF, 1'd0, 2'd1};
    ird_lut['h07a] = {UA_CALF, 1'd0, 2'd1};
    ird_lut['h07b] = {UA_CALF, 1'd0, 2'd1};
    ird_lut['h07c] = {UA_CALF, 1'd0, 2'd1};
    ird_lut['h07d] = {UA_CALF, 1'd0, 2'd1};
    ird_lut['h07e] = {UA_CALF, 1'd0, 2'd1};
    ird_lut['h07f] = {UA_CALF, 1'd0, 2'd1};
    ird_lut['h080] = {UA_CALT, 1'd0, 2'd0};
    ird_lut['h081] = {UA_CALT, 1'd0, 2'd0};
    ird_lut['h082] = {UA_CALT, 1'd0, 2'd0};
    ird_lut['h083] = {UA_CALT, 1'd0, 2'd0};
    ird_lut['h084] = {UA_CALT, 1'd0, 2'd0};
    ird_lut['h085] = {UA_CALT, 1'd0, 2'd0};
    ird_lut['h086] = {UA_CALT, 1'd0, 2'd0};
    ird_lut['h087] = {UA_CALT, 1'd0, 2'd0};
    ird_lut['h088] = {UA_CALT, 1'd0, 2'd0};
    ird_lut['h089] = {UA_CALT, 1'd0, 2'd0};
    ird_lut['h08a] = {UA_CALT, 1'd0, 2'd0};
    ird_lut['h08b] = {UA_CALT, 1'd0, 2'd0};
    ird_lut['h08c] = {UA_CALT, 1'd0, 2'd0};
    ird_lut['h08d] = {UA_CALT, 1'd0, 2'd0};
    ird_lut['h08e] = {UA_CALT, 1'd0, 2'd0};
    ird_lut['h08f] = {UA_CALT, 1'd0, 2'd0};
    ird_lut['h090] = {UA_CALT, 1'd0, 2'd0};
    ird_lut['h091] = {UA_CALT, 1'd0, 2'd0};
    ird_lut['h092] = {UA_CALT, 1'd0, 2'd0};
    ird_lut['h093] = {UA_CALT, 1'd0, 2'd0};
    ird_lut['h094] = {UA_CALT, 1'd0, 2'd0};
    ird_lut['h095] = {UA_CALT, 1'd0, 2'd0};
    ird_lut['h096] = {UA_CALT, 1'd0, 2'd0};
    ird_lut['h097] = {UA_CALT, 1'd0, 2'd0};
    ird_lut['h098] = {UA_CALT, 1'd0, 2'd0};
    ird_lut['h099] = {UA_CALT, 1'd0, 2'd0};
    ird_lut['h09a] = {UA_CALT, 1'd0, 2'd0};
    ird_lut['h09b] = {UA_CALT, 1'd0, 2'd0};
    ird_lut['h09c] = {UA_CALT, 1'd0, 2'd0};
    ird_lut['h09d] = {UA_CALT, 1'd0, 2'd0};
    ird_lut['h09e] = {UA_CALT, 1'd0, 2'd0};
    ird_lut['h09f] = {UA_CALT, 1'd0, 2'd0};
    ird_lut['h0a0] = {UA_CALT, 1'd0, 2'd0};
    ird_lut['h0a1] = {UA_CALT, 1'd0, 2'd0};
    ird_lut['h0a2] = {UA_CALT, 1'd0, 2'd0};
    ird_lut['h0a3] = {UA_CALT, 1'd0, 2'd0};
    ird_lut['h0a4] = {UA_CALT, 1'd0, 2'd0};
    ird_lut['h0a5] = {UA_CALT, 1'd0, 2'd0};
    ird_lut['h0a6] = {UA_CALT, 1'd0, 2'd0};
    ird_lut['h0a7] = {UA_CALT, 1'd0, 2'd0};
    ird_lut['h0a8] = {UA_CALT, 1'd0, 2'd0};
    ird_lut['h0a9] = {UA_CALT, 1'd0, 2'd0};
    ird_lut['h0aa] = {UA_CALT, 1'd0, 2'd0};
    ird_lut['h0ab] = {UA_CALT, 1'd0, 2'd0};
    ird_lut['h0ac] = {UA_CALT, 1'd0, 2'd0};
    ird_lut['h0ad] = {UA_CALT, 1'd0, 2'd0};
    ird_lut['h0ae] = {UA_CALT, 1'd0, 2'd0};
    ird_lut['h0af] = {UA_CALT, 1'd0, 2'd0};
    ird_lut['h0b0] = {UA_CALT, 1'd0, 2'd0};
    ird_lut['h0b1] = {UA_CALT, 1'd0, 2'd0};
    ird_lut['h0b2] = {UA_CALT, 1'd0, 2'd0};
    ird_lut['h0b3] = {UA_CALT, 1'd0, 2'd0};
    ird_lut['h0b4] = {UA_CALT, 1'd0, 2'd0};
    ird_lut['h0b5] = {UA_CALT, 1'd0, 2'd0};
    ird_lut['h0b6] = {UA_CALT, 1'd0, 2'd0};
    ird_lut['h0b7] = {UA_CALT, 1'd0, 2'd0};
    ird_lut['h0b8] = {UA_CALT, 1'd0, 2'd0};
    ird_lut['h0b9] = {UA_CALT, 1'd0, 2'd0};
    ird_lut['h0ba] = {UA_CALT, 1'd0, 2'd0};
    ird_lut['h0bb] = {UA_CALT, 1'd0, 2'd0};
    ird_lut['h0bc] = {UA_CALT, 1'd0, 2'd0};
    ird_lut['h0bd] = {UA_CALT, 1'd0, 2'd0};
    ird_lut['h0be] = {UA_CALT, 1'd0, 2'd0};
    ird_lut['h0bf] = {UA_CALT, 1'd0, 2'd0};
    ird_lut['h072] = {UA_INT, 1'd0, 2'd0};
    ird_lut['h008] = {UA_RET, 1'd0, 2'd0};
    ird_lut['h062] = {UA_RETI, 1'd0, 2'd0};
    ird_lut['h058] = {UA_BIT, 1'd0, 2'd1};
    ird_lut['h059] = {UA_BIT, 1'd0, 2'd1};
    ird_lut['h05a] = {UA_BIT, 1'd0, 2'd1};
    ird_lut['h05b] = {UA_BIT, 1'd0, 2'd1};
    ird_lut['h05c] = {UA_BIT, 1'd0, 2'd1};
    ird_lut['h05d] = {UA_BIT, 1'd0, 2'd1};
    ird_lut['h05e] = {UA_BIT, 1'd0, 2'd1};
    ird_lut['h05f] = {UA_BIT, 1'd0, 2'd1};
    ird_lut['h000] = {UA_IDLE, 1'd1, 2'd0};
    ird_lut['h019] = {UA_STM, 1'd1, 2'd0};
    ird_lut['h130] = {UA_RLL_A_, 1'd1, 2'd0};
    ird_lut['h131] = {UA_RLR_A_, 1'd1, 2'd0};
    ird_lut['h132] = {UA_RLL_C_, 1'd1, 2'd0};
    ird_lut['h133] = {UA_RLR_C_, 1'd1, 2'd0};
    ird_lut['h134] = {UA_SLL_A_, 1'd1, 2'd0};
    ird_lut['h135] = {UA_SLR_A_, 1'd1, 2'd0};
    ird_lut['h136] = {UA_SLL_C_, 1'd1, 2'd0};
    ird_lut['h137] = {UA_SLR_C_, 1'd1, 2'd0};
    ird_lut['h10e] = {UA_PUSH_VA, 1'd0, 2'd0};
    ird_lut['h10f] = {UA_POP_VA, 1'd0, 2'd0};
    ird_lut['h11e] = {UA_PUSH_BC, 1'd0, 2'd0};
    ird_lut['h11f] = {UA_POP_BC, 1'd0, 2'd0};
    ird_lut['h12e] = {UA_PUSH_DE, 1'd0, 2'd0};
    ird_lut['h12f] = {UA_POP_DE, 1'd0, 2'd0};
    ird_lut['h13e] = {UA_PUSH_HL, 1'd0, 2'd0};
    ird_lut['h13f] = {UA_POP_HL, 1'd0, 2'd0};
    ird_lut['h100] = {UA_SKIP_I, 1'd1, 2'd0};
    ird_lut['h101] = {UA_SKIP_I, 1'd1, 2'd0};
    ird_lut['h102] = {UA_SKIP_I, 1'd1, 2'd0};
    ird_lut['h103] = {UA_SKIP_I, 1'd1, 2'd0};
    ird_lut['h104] = {UA_SKIP_I, 1'd1, 2'd0};
    ird_lut['h10a] = {UA_SKIP_C, 1'd1, 2'd0};
    ird_lut['h110] = {UA_SKIP_NI, 1'd1, 2'd0};
    ird_lut['h111] = {UA_SKIP_NI, 1'd1, 2'd0};
    ird_lut['h112] = {UA_SKIP_NI, 1'd1, 2'd0};
    ird_lut['h113] = {UA_SKIP_NI, 1'd1, 2'd0};
    ird_lut['h114] = {UA_SKIP_NI, 1'd1, 2'd0};
    ird_lut['h11a] = {UA_SKIP_NC, 1'd1, 2'd0};
    ird_lut['h120] = {UA_EI, 1'd1, 2'd0};
    ird_lut['h124] = {UA_DI, 1'd1, 2'd0};
    ird_lut['h2c0] = {UA_MOV_A_SPR_IR3, 1'd1, 2'd0};
    ird_lut['h2c1] = {UA_MOV_A_SPR_IR3, 1'd1, 2'd0};
    ird_lut['h2c2] = {UA_MOV_A_SPR_IR3, 1'd1, 2'd0};
    ird_lut['h2c3] = {UA_MOV_A_SPR_IR3, 1'd1, 2'd0};
    ird_lut['h2c4] = {UA_MOV_A_SPR_IR3, 1'd1, 2'd0};
    ird_lut['h2c5] = {UA_MOV_A_SPR_IR3, 1'd1, 2'd0};
    ird_lut['h2c6] = {UA_MOV_A_SPR_IR3, 1'd1, 2'd0};
    ird_lut['h2c7] = {UA_MOV_A_SPR_IR3, 1'd1, 2'd0};
    ird_lut['h2c8] = {UA_MOV_A_SPR_IR3, 1'd1, 2'd0};
    ird_lut['h2c9] = {UA_MOV_A_SPR_IR3, 1'd1, 2'd0};
    ird_lut['h3c0] = {UA_MOV_SPR_IR3_A, 1'd1, 2'd0};
    ird_lut['h3c1] = {UA_MOV_SPR_IR3_A, 1'd1, 2'd0};
    ird_lut['h3c2] = {UA_MOV_SPR_IR3_A, 1'd1, 2'd0};
    ird_lut['h3c3] = {UA_MOV_SPR_IR3_A, 1'd1, 2'd0};
    ird_lut['h3c4] = {UA_MOV_SPR_IR3_A, 1'd1, 2'd0};
    ird_lut['h3c5] = {UA_MOV_SPR_IR3_A, 1'd1, 2'd0};
    ird_lut['h3c6] = {UA_MOV_SPR_IR3_A, 1'd1, 2'd0};
    ird_lut['h3c7] = {UA_MOV_SPR_IR3_A, 1'd1, 2'd0};
    ird_lut['h3c8] = {UA_MOV_SPR_IR3_A, 1'd1, 2'd0};
    ird_lut['h3c9] = {UA_MOV_SPR_IR3_A, 1'd1, 2'd0};
    ird_lut['h420] = {UA_ADDNC_RF_IR210_A, 1'd1, 2'd0};
    ird_lut['h421] = {UA_ADDNC_RF_IR210_A, 1'd1, 2'd0};
    ird_lut['h422] = {UA_ADDNC_RF_IR210_A, 1'd1, 2'd0};
    ird_lut['h423] = {UA_ADDNC_RF_IR210_A, 1'd1, 2'd0};
    ird_lut['h424] = {UA_ADDNC_RF_IR210_A, 1'd1, 2'd0};
    ird_lut['h425] = {UA_ADDNC_RF_IR210_A, 1'd1, 2'd0};
    ird_lut['h426] = {UA_ADDNC_RF_IR210_A, 1'd1, 2'd0};
    ird_lut['h427] = {UA_ADDNC_RF_IR210_A, 1'd1, 2'd0};
    ird_lut['h430] = {UA_SUBNB_RF_IR210_A, 1'd1, 2'd0};
    ird_lut['h431] = {UA_SUBNB_RF_IR210_A, 1'd1, 2'd0};
    ird_lut['h432] = {UA_SUBNB_RF_IR210_A, 1'd1, 2'd0};
    ird_lut['h433] = {UA_SUBNB_RF_IR210_A, 1'd1, 2'd0};
    ird_lut['h434] = {UA_SUBNB_RF_IR210_A, 1'd1, 2'd0};
    ird_lut['h435] = {UA_SUBNB_RF_IR210_A, 1'd1, 2'd0};
    ird_lut['h436] = {UA_SUBNB_RF_IR210_A, 1'd1, 2'd0};
    ird_lut['h437] = {UA_SUBNB_RF_IR210_A, 1'd1, 2'd0};
    ird_lut['h440] = {UA_ADD_RF_IR210_A, 1'd1, 2'd0};
    ird_lut['h441] = {UA_ADD_RF_IR210_A, 1'd1, 2'd0};
    ird_lut['h442] = {UA_ADD_RF_IR210_A, 1'd1, 2'd0};
    ird_lut['h443] = {UA_ADD_RF_IR210_A, 1'd1, 2'd0};
    ird_lut['h444] = {UA_ADD_RF_IR210_A, 1'd1, 2'd0};
    ird_lut['h445] = {UA_ADD_RF_IR210_A, 1'd1, 2'd0};
    ird_lut['h446] = {UA_ADD_RF_IR210_A, 1'd1, 2'd0};
    ird_lut['h447] = {UA_ADD_RF_IR210_A, 1'd1, 2'd0};
    ird_lut['h450] = {UA_ADC_RF_IR210_A, 1'd1, 2'd0};
    ird_lut['h451] = {UA_ADC_RF_IR210_A, 1'd1, 2'd0};
    ird_lut['h452] = {UA_ADC_RF_IR210_A, 1'd1, 2'd0};
    ird_lut['h453] = {UA_ADC_RF_IR210_A, 1'd1, 2'd0};
    ird_lut['h454] = {UA_ADC_RF_IR210_A, 1'd1, 2'd0};
    ird_lut['h455] = {UA_ADC_RF_IR210_A, 1'd1, 2'd0};
    ird_lut['h456] = {UA_ADC_RF_IR210_A, 1'd1, 2'd0};
    ird_lut['h457] = {UA_ADC_RF_IR210_A, 1'd1, 2'd0};
    ird_lut['h460] = {UA_SUB_RF_IR210_A, 1'd1, 2'd0};
    ird_lut['h461] = {UA_SUB_RF_IR210_A, 1'd1, 2'd0};
    ird_lut['h462] = {UA_SUB_RF_IR210_A, 1'd1, 2'd0};
    ird_lut['h463] = {UA_SUB_RF_IR210_A, 1'd1, 2'd0};
    ird_lut['h464] = {UA_SUB_RF_IR210_A, 1'd1, 2'd0};
    ird_lut['h465] = {UA_SUB_RF_IR210_A, 1'd1, 2'd0};
    ird_lut['h466] = {UA_SUB_RF_IR210_A, 1'd1, 2'd0};
    ird_lut['h467] = {UA_SUB_RF_IR210_A, 1'd1, 2'd0};
    ird_lut['h470] = {UA_SBB_RF_IR210_A, 1'd1, 2'd0};
    ird_lut['h471] = {UA_SBB_RF_IR210_A, 1'd1, 2'd0};
    ird_lut['h472] = {UA_SBB_RF_IR210_A, 1'd1, 2'd0};
    ird_lut['h473] = {UA_SBB_RF_IR210_A, 1'd1, 2'd0};
    ird_lut['h474] = {UA_SBB_RF_IR210_A, 1'd1, 2'd0};
    ird_lut['h475] = {UA_SBB_RF_IR210_A, 1'd1, 2'd0};
    ird_lut['h476] = {UA_SBB_RF_IR210_A, 1'd1, 2'd0};
    ird_lut['h477] = {UA_SBB_RF_IR210_A, 1'd1, 2'd0};
    ird_lut['h4b0] = {UA_SUBNB_A_RF_IR210, 1'd1, 2'd0};
    ird_lut['h4b1] = {UA_SUBNB_A_RF_IR210, 1'd1, 2'd0};
    ird_lut['h4b2] = {UA_SUBNB_A_RF_IR210, 1'd1, 2'd0};
    ird_lut['h4b3] = {UA_SUBNB_A_RF_IR210, 1'd1, 2'd0};
    ird_lut['h4b4] = {UA_SUBNB_A_RF_IR210, 1'd1, 2'd0};
    ird_lut['h4b5] = {UA_SUBNB_A_RF_IR210, 1'd1, 2'd0};
    ird_lut['h4b6] = {UA_SUBNB_A_RF_IR210, 1'd1, 2'd0};
    ird_lut['h4b7] = {UA_SUBNB_A_RF_IR210, 1'd1, 2'd0};
    ird_lut['h4c0] = {UA_ADD_A_RF_IR210, 1'd1, 2'd0};
    ird_lut['h4c1] = {UA_ADD_A_RF_IR210, 1'd1, 2'd0};
    ird_lut['h4c2] = {UA_ADD_A_RF_IR210, 1'd1, 2'd0};
    ird_lut['h4c3] = {UA_ADD_A_RF_IR210, 1'd1, 2'd0};
    ird_lut['h4c4] = {UA_ADD_A_RF_IR210, 1'd1, 2'd0};
    ird_lut['h4c5] = {UA_ADD_A_RF_IR210, 1'd1, 2'd0};
    ird_lut['h4c6] = {UA_ADD_A_RF_IR210, 1'd1, 2'd0};
    ird_lut['h4c7] = {UA_ADD_A_RF_IR210, 1'd1, 2'd0};
    ird_lut['h4d0] = {UA_ADC_A_RF_IR210, 1'd1, 2'd0};
    ird_lut['h4d1] = {UA_ADC_A_RF_IR210, 1'd1, 2'd0};
    ird_lut['h4d2] = {UA_ADC_A_RF_IR210, 1'd1, 2'd0};
    ird_lut['h4d3] = {UA_ADC_A_RF_IR210, 1'd1, 2'd0};
    ird_lut['h4d4] = {UA_ADC_A_RF_IR210, 1'd1, 2'd0};
    ird_lut['h4d5] = {UA_ADC_A_RF_IR210, 1'd1, 2'd0};
    ird_lut['h4d6] = {UA_ADC_A_RF_IR210, 1'd1, 2'd0};
    ird_lut['h4d7] = {UA_ADC_A_RF_IR210, 1'd1, 2'd0};
    ird_lut['h4e0] = {UA_SUB_A_RF_IR210, 1'd1, 2'd0};
    ird_lut['h4e1] = {UA_SUB_A_RF_IR210, 1'd1, 2'd0};
    ird_lut['h4e2] = {UA_SUB_A_RF_IR210, 1'd1, 2'd0};
    ird_lut['h4e3] = {UA_SUB_A_RF_IR210, 1'd1, 2'd0};
    ird_lut['h4e4] = {UA_SUB_A_RF_IR210, 1'd1, 2'd0};
    ird_lut['h4e5] = {UA_SUB_A_RF_IR210, 1'd1, 2'd0};
    ird_lut['h4e6] = {UA_SUB_A_RF_IR210, 1'd1, 2'd0};
    ird_lut['h4e7] = {UA_SUB_A_RF_IR210, 1'd1, 2'd0};
    ird_lut['h4f0] = {UA_SBB_A_RF_IR210, 1'd1, 2'd0};
    ird_lut['h4f1] = {UA_SBB_A_RF_IR210, 1'd1, 2'd0};
    ird_lut['h4f2] = {UA_SBB_A_RF_IR210, 1'd1, 2'd0};
    ird_lut['h4f3] = {UA_SBB_A_RF_IR210, 1'd1, 2'd0};
    ird_lut['h4f4] = {UA_SBB_A_RF_IR210, 1'd1, 2'd0};
    ird_lut['h4f5] = {UA_SBB_A_RF_IR210, 1'd1, 2'd0};
    ird_lut['h4f6] = {UA_SBB_A_RF_IR210, 1'd1, 2'd0};
    ird_lut['h4f7] = {UA_SBB_A_RF_IR210, 1'd1, 2'd0};
    ird_lut['h520] = {UA_ADDNC_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h521] = {UA_ADDNC_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h522] = {UA_ADDNC_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h523] = {UA_ADDNC_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h524] = {UA_ADDNC_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h525] = {UA_ADDNC_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h526] = {UA_ADDNC_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h527] = {UA_ADDNC_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h530] = {UA_SUBNB_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h531] = {UA_SUBNB_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h532] = {UA_SUBNB_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h533] = {UA_SUBNB_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h534] = {UA_SUBNB_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h535] = {UA_SUBNB_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h536] = {UA_SUBNB_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h537] = {UA_SUBNB_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h540] = {UA_ADD_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h541] = {UA_ADD_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h542] = {UA_ADD_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h543] = {UA_ADD_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h544] = {UA_ADD_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h545] = {UA_ADD_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h546] = {UA_ADD_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h547] = {UA_ADD_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h550] = {UA_ADC_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h551] = {UA_ADC_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h552] = {UA_ADC_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h553] = {UA_ADC_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h554] = {UA_ADC_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h555] = {UA_ADC_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h556] = {UA_ADC_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h557] = {UA_ADC_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h558] = {UA_OFF_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h559] = {UA_OFF_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h55a] = {UA_OFF_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h55b] = {UA_OFF_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h55c] = {UA_OFF_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h55d] = {UA_OFF_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h55e] = {UA_OFF_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h55f] = {UA_OFF_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h560] = {UA_SUB_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h561] = {UA_SUB_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h562] = {UA_SUB_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h563] = {UA_SUB_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h564] = {UA_SUB_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h565] = {UA_SUB_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h566] = {UA_SUB_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h567] = {UA_SUB_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h570] = {UA_SBB_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h571] = {UA_SBB_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h572] = {UA_SBB_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h573] = {UA_SBB_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h574] = {UA_SBB_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h575] = {UA_SBB_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h576] = {UA_SBB_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h577] = {UA_SBB_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h588] = {UA_AND_SPR_IR2_IMM, 1'd0, 2'd1};
    ird_lut['h589] = {UA_AND_SPR_IR2_IMM, 1'd0, 2'd1};
    ird_lut['h58a] = {UA_AND_SPR_IR2_IMM, 1'd0, 2'd1};
    ird_lut['h58b] = {UA_AND_SPR_IR2_IMM, 1'd0, 2'd1};
    ird_lut['h58c] = {UA_AND_SPR_IR2_IMM, 1'd0, 2'd1};
    ird_lut['h58d] = {UA_AND_SPR_IR2_IMM, 1'd0, 2'd1};
    ird_lut['h58e] = {UA_AND_SPR_IR2_IMM, 1'd0, 2'd1};
    ird_lut['h58f] = {UA_AND_SPR_IR2_IMM, 1'd0, 2'd1};
    ird_lut['h590] = {UA_XOR_SPR_IR2_IMM, 1'd0, 2'd1};
    ird_lut['h591] = {UA_XOR_SPR_IR2_IMM, 1'd0, 2'd1};
    ird_lut['h592] = {UA_XOR_SPR_IR2_IMM, 1'd0, 2'd1};
    ird_lut['h593] = {UA_XOR_SPR_IR2_IMM, 1'd0, 2'd1};
    ird_lut['h594] = {UA_XOR_SPR_IR2_IMM, 1'd0, 2'd1};
    ird_lut['h595] = {UA_XOR_SPR_IR2_IMM, 1'd0, 2'd1};
    ird_lut['h596] = {UA_XOR_SPR_IR2_IMM, 1'd0, 2'd1};
    ird_lut['h597] = {UA_XOR_SPR_IR2_IMM, 1'd0, 2'd1};
    ird_lut['h598] = {UA_OR_SPR_IR2_IMM, 1'd0, 2'd1};
    ird_lut['h599] = {UA_OR_SPR_IR2_IMM, 1'd0, 2'd1};
    ird_lut['h59a] = {UA_OR_SPR_IR2_IMM, 1'd0, 2'd1};
    ird_lut['h59b] = {UA_OR_SPR_IR2_IMM, 1'd0, 2'd1};
    ird_lut['h59c] = {UA_OR_SPR_IR2_IMM, 1'd0, 2'd1};
    ird_lut['h59d] = {UA_OR_SPR_IR2_IMM, 1'd0, 2'd1};
    ird_lut['h59e] = {UA_OR_SPR_IR2_IMM, 1'd0, 2'd1};
    ird_lut['h59f] = {UA_OR_SPR_IR2_IMM, 1'd0, 2'd1};
    ird_lut['h548] = {UA_ON_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h549] = {UA_ON_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h54a] = {UA_ON_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h54b] = {UA_ON_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h54c] = {UA_ON_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h54d] = {UA_ON_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h54e] = {UA_ON_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h54f] = {UA_ON_RF_IR210_IMM, 1'd0, 2'd1};
    ird_lut['h5c8] = {UA_ON_SPR_IR2_IMM, 1'd0, 2'd1};
    ird_lut['h5c9] = {UA_ON_SPR_IR2_IMM, 1'd0, 2'd1};
    ird_lut['h5ca] = {UA_ON_SPR_IR2_IMM, 1'd0, 2'd1};
    ird_lut['h5cb] = {UA_ON_SPR_IR2_IMM, 1'd0, 2'd1};
    ird_lut['h5cc] = {UA_ON_SPR_IR2_IMM, 1'd0, 2'd1};
    ird_lut['h5cd] = {UA_ON_SPR_IR2_IMM, 1'd0, 2'd1};
    ird_lut['h5ce] = {UA_ON_SPR_IR2_IMM, 1'd0, 2'd1};
    ird_lut['h5cf] = {UA_ON_SPR_IR2_IMM, 1'd0, 2'd1};
    ird_lut['h5d8] = {UA_OFF_SPR_IR2_IMM, 1'd0, 2'd1};
    ird_lut['h5d9] = {UA_OFF_SPR_IR2_IMM, 1'd0, 2'd1};
    ird_lut['h5da] = {UA_OFF_SPR_IR2_IMM, 1'd0, 2'd1};
    ird_lut['h5db] = {UA_OFF_SPR_IR2_IMM, 1'd0, 2'd1};
    ird_lut['h5dc] = {UA_OFF_SPR_IR2_IMM, 1'd0, 2'd1};
    ird_lut['h5dd] = {UA_OFF_SPR_IR2_IMM, 1'd0, 2'd1};
    ird_lut['h5de] = {UA_OFF_SPR_IR2_IMM, 1'd0, 2'd1};
    ird_lut['h5df] = {UA_OFF_SPR_IR2_IMM, 1'd0, 2'd1};
    ird_lut['h668] = {UA_LD_IR210_ABS, 1'd0, 2'd2};
    ird_lut['h669] = {UA_LD_IR210_ABS, 1'd0, 2'd2};
    ird_lut['h66a] = {UA_LD_IR210_ABS, 1'd0, 2'd2};
    ird_lut['h66b] = {UA_LD_IR210_ABS, 1'd0, 2'd2};
    ird_lut['h66c] = {UA_LD_IR210_ABS, 1'd0, 2'd2};
    ird_lut['h66d] = {UA_LD_IR210_ABS, 1'd0, 2'd2};
    ird_lut['h66e] = {UA_LD_IR210_ABS, 1'd0, 2'd2};
    ird_lut['h66f] = {UA_LD_IR210_ABS, 1'd0, 2'd2};
    ird_lut['h678] = {UA_ST_IR210_ABS, 1'd0, 2'd2};
    ird_lut['h679] = {UA_ST_IR210_ABS, 1'd0, 2'd2};
    ird_lut['h67a] = {UA_ST_IR210_ABS, 1'd0, 2'd2};
    ird_lut['h67b] = {UA_ST_IR210_ABS, 1'd0, 2'd2};
    ird_lut['h67c] = {UA_ST_IR210_ABS, 1'd0, 2'd2};
    ird_lut['h67d] = {UA_ST_IR210_ABS, 1'd0, 2'd2};
    ird_lut['h67e] = {UA_ST_IR210_ABS, 1'd0, 2'd2};
    ird_lut['h67f] = {UA_ST_IR210_ABS, 1'd0, 2'd2};
    ird_lut['h6c1] = {UA_ADD, 1'd0, 2'd0};
    ird_lut['h6c2] = {UA_ADD, 1'd0, 2'd0};
    ird_lut['h6c3] = {UA_ADD, 1'd0, 2'd0};
    ird_lut['h6c4] = {UA_ADD, 1'd0, 2'd0};
    ird_lut['h6c5] = {UA_ADD, 1'd0, 2'd0};
    ird_lut['h6c6] = {UA_ADD, 1'd0, 2'd0};
    ird_lut['h6c7] = {UA_ADD, 1'd0, 2'd0};
    ird_lut['h6e1] = {UA_SUB, 1'd0, 2'd0};
    ird_lut['h6e2] = {UA_SUB, 1'd0, 2'd0};
    ird_lut['h6e3] = {UA_SUB, 1'd0, 2'd0};
    ird_lut['h6e4] = {UA_SUB, 1'd0, 2'd0};
    ird_lut['h6e5] = {UA_SUB, 1'd0, 2'd0};
    ird_lut['h6e6] = {UA_SUB, 1'd0, 2'd0};
    ird_lut['h6e7] = {UA_SUB, 1'd0, 2'd0};
    ird_lut['h7c0] = {UA_ADD_A_WA, 1'd0, 2'd1};
    ird_lut['h788] = {UA_AND_A_WA, 1'd0, 2'd1};
    ird_lut['h798] = {UA_OR_A_WA, 1'd0, 2'd1};
