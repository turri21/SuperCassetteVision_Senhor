typedef enum reg [9:0]
{
    UA_IDLE,
    UA_SKIP_OP2,
    UA__2,
    UA__3,
    UA_SKIP_OP1,
    UA__5,
    UA__6,
    UA_MOV_A_RF_IR210,
    UA__8,
    UA__9,
    UA_MOV_RF_IR210_A,
    UA__B,
    UA__C,
    UA_MOV_RF_IR210_IMM,
    UA__E,
    UA__F,
    UA_LD_A_WA,
    UA__11,
    UA__12,
    UA__13,
    UA__14,
    UA__15,
    UA_LDX_SP_IMM,
    UA__17,
    UA__18,
    UA__19,
    UA__1A,
    UA__1B,
    UA_LDX_BC_IMM,
    UA__1D,
    UA__1E,
    UA__1F,
    UA__20,
    UA__21,
    UA_LDX_DE_IMM,
    UA__23,
    UA__24,
    UA__25,
    UA__26,
    UA__27,
    UA_LDX_HL_IMM,
    UA__29,
    UA__2A,
    UA__2B,
    UA__2C,
    UA__2D,
    UA_LDAX,
    UA__2F,
    UA__30,
    UA_STX_A,
    UA__32,
    UA__33,
    UA_STX_RF_W,
    UA__35,
    UA__36,
    UA__37,
    UA__38,
    UA__39,
    UA_STW_A,
    UA__3B,
    UA__3C,
    UA__3D,
    UA__3E,
    UA__3F,
    UA_STW_IMM,
    UA__41,
    UA__42,
    UA__43,
    UA__44,
    UA__45,
    UA__46,
    UA__47,
    UA__48,
    UA_TABLE,
    UA__4A,
    UA__4B,
    UA__4C,
    UA__4D,
    UA__4E,
    UA__4F,
    UA__50,
    UA__51,
    UA__52,
    UA__53,
    UA__54,
    UA__55,
    UA__56,
    UA__57,
    UA_BLOCK,
    UA__59,
    UA__5A,
    UA__5B,
    UA__5C,
    UA__5D,
    UA__5E,
    UA__5F,
    UA__60,
    UA_AND_WA_IMM,
    UA__62,
    UA__63,
    UA__64,
    UA__65,
    UA__66,
    UA__67,
    UA__68,
    UA__69,
    UA__6A,
    UA__6B,
    UA__6C,
    UA_OR_WA_IMM,
    UA__6E,
    UA__6F,
    UA__70,
    UA__71,
    UA__72,
    UA__73,
    UA__74,
    UA__75,
    UA__76,
    UA__77,
    UA__78,
    UA_AND_A_IMM,
    UA__7A,
    UA__7B,
    UA__7C,
    UA_XOR_A_IMM,
    UA__7E,
    UA__7F,
    UA__80,
    UA_OR_A_IMM,
    UA__82,
    UA__83,
    UA__84,
    UA_CMPBNB_WA_IMM,
    UA__86,
    UA__87,
    UA__88,
    UA__89,
    UA__8A,
    UA__8B,
    UA__8C,
    UA__8D,
    UA__8E,
    UA_CMPB_WA_IMM,
    UA__90,
    UA__91,
    UA__92,
    UA__93,
    UA__94,
    UA__95,
    UA__96,
    UA__97,
    UA__98,
    UA_BITNZ_WA_IMM,
    UA__9A,
    UA__9B,
    UA__9C,
    UA__9D,
    UA__9E,
    UA__9F,
    UA__A0,
    UA__A1,
    UA__A2,
    UA_BITZ_WA_IMM,
    UA__A4,
    UA__A5,
    UA__A6,
    UA__A7,
    UA__A8,
    UA__A9,
    UA__AA,
    UA__AB,
    UA__AC,
    UA_CMPNZ_WA_IMM,
    UA__AE,
    UA__AF,
    UA__B0,
    UA__B1,
    UA__B2,
    UA__B3,
    UA__B4,
    UA__B5,
    UA__B6,
    UA_CMPZ_WA_IMM,
    UA__B8,
    UA__B9,
    UA__BA,
    UA__BB,
    UA__BC,
    UA__BD,
    UA__BE,
    UA__BF,
    UA__C0,
    UA_CMPBNB_A_IMM,
    UA__C2,
    UA__C3,
    UA__C4,
    UA_CMPB_A_IMM,
    UA__C6,
    UA__C7,
    UA__C8,
    UA_BITNZ_A_IMM,
    UA__CA,
    UA__CB,
    UA__CC,
    UA_BITZ_A_IMM,
    UA__CE,
    UA__CF,
    UA__D0,
    UA_CMPNZ_A_IMM,
    UA__D2,
    UA__D3,
    UA__D4,
    UA_CMPZ_A_IMM,
    UA__D6,
    UA__D7,
    UA__D8,
    UA_ADDNC_A_IMM,
    UA__DA,
    UA__DB,
    UA__DC,
    UA_SUBNB_A_IMM,
    UA__DE,
    UA__DF,
    UA__E0,
    UA_ADD_A_IMM,
    UA__E2,
    UA__E3,
    UA__E4,
    UA_ADC_A_IMM,
    UA__E6,
    UA__E7,
    UA__E8,
    UA_SUB_A_IMM,
    UA__EA,
    UA__EB,
    UA__EC,
    UA_SBB_A_IMM,
    UA__EE,
    UA__EF,
    UA__F0,
    UA_INCR_WA,
    UA__F2,
    UA__F3,
    UA__F4,
    UA__F5,
    UA__F6,
    UA__F7,
    UA__F8,
    UA__F9,
    UA_DECR_WA,
    UA__FB,
    UA__FC,
    UA__FD,
    UA__FE,
    UA__FF,
    UA__100,
    UA__101,
    UA__102,
    UA_INCR_RF_IR210,
    UA__104,
    UA_DECR_RF_IR210,
    UA__106,
    UA_INC_SP,
    UA__108,
    UA__109,
    UA_INC_BC,
    UA__10B,
    UA__10C,
    UA_INC_DE,
    UA__10E,
    UA__10F,
    UA_INC_HL,
    UA__111,
    UA__112,
    UA_DEC_SP,
    UA__114,
    UA__115,
    UA_DEC_BC,
    UA__117,
    UA__118,
    UA_DEC_DE,
    UA__11A,
    UA__11B,
    UA_DEC_HL,
    UA__11D,
    UA__11E,
    UA_DAA,
    UA__120,
    UA_JR,
    UA__122,
    UA__123,
    UA__124,
    UA__125,
    UA__126,
    UA__127,
    UA__128,
    UA__129,
    UA_JRE_P,
    UA__12B,
    UA__12C,
    UA__12D,
    UA__12E,
    UA__12F,
    UA__130,
    UA__131,
    UA__132,
    UA_JRE_N,
    UA__134,
    UA__135,
    UA__136,
    UA__137,
    UA__138,
    UA__139,
    UA__13A,
    UA__13B,
    UA_JMP,
    UA__13D,
    UA__13E,
    UA__13F,
    UA__140,
    UA__141,
    UA_JB,
    UA_CALL,
    UA__144,
    UA__145,
    UA__146,
    UA__147,
    UA__148,
    UA__149,
    UA__14A,
    UA__14B,
    UA__14C,
    UA__14D,
    UA__14E,
    UA_CALB,
    UA__150,
    UA__151,
    UA__152,
    UA__153,
    UA__154,
    UA__155,
    UA__156,
    UA__157,
    UA_CALF,
    UA__159,
    UA__15A,
    UA__15B,
    UA__15C,
    UA__15D,
    UA__15E,
    UA__15F,
    UA__160,
    UA__161,
    UA__162,
    UA__163,
    UA_CALT,
    UA__165,
    UA__166,
    UA__167,
    UA__168,
    UA__169,
    UA__16A,
    UA__16B,
    UA__16C,
    UA__16D,
    UA__16E,
    UA__16F,
    UA__170,
    UA__171,
    UA__172,
    UA_INT,
    UA__174,
    UA__175,
    UA__176,
    UA__177,
    UA__178,
    UA__179,
    UA__17A,
    UA__17B,
    UA__17C,
    UA__17D,
    UA__17E,
    UA__17F,
    UA__180,
    UA__181,
    UA__182,
    UA__183,
    UA__184,
    UA_RET,
    UA__186,
    UA__187,
    UA__188,
    UA__189,
    UA__18A,
    UA_RETS,
    UA__18C,
    UA__18D,
    UA__18E,
    UA__18F,
    UA__190,
    UA_RETI,
    UA__192,
    UA__193,
    UA__194,
    UA__195,
    UA__196,
    UA__197,
    UA__198,
    UA__199,
    UA_BIT,
    UA__19B,
    UA__19C,
    UA__19D,
    UA__19E,
    UA__19F,
    UA__1A0,
    UA_STM,
    UA_RLL_A_,
    UA__1A3,
    UA__1A4,
    UA_RLR_A_,
    UA__1A6,
    UA__1A7,
    UA_RLL_C_,
    UA__1A9,
    UA__1AA,
    UA_RLR_C_,
    UA__1AC,
    UA__1AD,
    UA_SLL_A_,
    UA__1AF,
    UA__1B0,
    UA_SLR_A_,
    UA__1B2,
    UA__1B3,
    UA_SLL_C_,
    UA__1B5,
    UA__1B6,
    UA_SLR_C_,
    UA__1B8,
    UA__1B9,
    UA_PUSH_VA,
    UA__1BB,
    UA__1BC,
    UA__1BD,
    UA__1BE,
    UA__1BF,
    UA__1C0,
    UA__1C1,
    UA__1C2,
    UA_POP_VA,
    UA__1C4,
    UA__1C5,
    UA__1C6,
    UA__1C7,
    UA__1C8,
    UA_PUSH_BC,
    UA__1CA,
    UA__1CB,
    UA__1CC,
    UA__1CD,
    UA__1CE,
    UA__1CF,
    UA__1D0,
    UA__1D1,
    UA_POP_BC,
    UA__1D3,
    UA__1D4,
    UA__1D5,
    UA__1D6,
    UA__1D7,
    UA_PUSH_DE,
    UA__1D9,
    UA__1DA,
    UA__1DB,
    UA__1DC,
    UA__1DD,
    UA__1DE,
    UA__1DF,
    UA__1E0,
    UA_POP_DE,
    UA__1E2,
    UA__1E3,
    UA__1E4,
    UA__1E5,
    UA__1E6,
    UA_PUSH_HL,
    UA__1E8,
    UA__1E9,
    UA__1EA,
    UA__1EB,
    UA__1EC,
    UA__1ED,
    UA__1EE,
    UA__1EF,
    UA_POP_HL,
    UA__1F1,
    UA__1F2,
    UA__1F3,
    UA__1F4,
    UA__1F5,
    UA_SKIP_I,
    UA_SKIP_PSW_C,
    UA_SKIP_PSW_Z,
    UA_SKIP_NI,
    UA_SKIP_PSW_NC,
    UA_SKIP_PSW_NZ,
    UA_EI,
    UA_DI,
    UA_CLC,
    UA_STC,
    UA_RLD,
    UA__201,
    UA__202,
    UA__203,
    UA__204,
    UA__205,
    UA__206,
    UA__207,
    UA__208,
    UA__209,
    UA_RRD,
    UA__20B,
    UA__20C,
    UA__20D,
    UA__20E,
    UA__20F,
    UA__210,
    UA__211,
    UA__212,
    UA__213,
    UA_MOV_A_SPR_IR3,
    UA__215,
    UA__216,
    UA_MOV_SPR_IR3_A,
    UA__218,
    UA__219,
    UA_ADDNC_RF_IR210_A,
    UA__21B,
    UA__21C,
    UA_SUBNB_RF_IR210_A,
    UA__21E,
    UA__21F,
    UA_ADD_RF_IR210_A,
    UA__221,
    UA__222,
    UA_ADC_RF_IR210_A,
    UA__224,
    UA__225,
    UA_SUB_RF_IR210_A,
    UA__227,
    UA__228,
    UA_SBB_RF_IR210_A,
    UA__22A,
    UA__22B,
    UA_ADDNC_A_RF_IR210,
    UA__22D,
    UA__22E,
    UA_SUBNB_A_RF_IR210,
    UA__230,
    UA__231,
    UA_ADD_A_RF_IR210,
    UA__233,
    UA__234,
    UA_ADC_A_RF_IR210,
    UA__236,
    UA__237,
    UA_SUB_A_RF_IR210,
    UA__239,
    UA__23A,
    UA_SBB_A_RF_IR210,
    UA__23C,
    UA__23D,
    UA_AND_RF_IR210_A,
    UA__23F,
    UA__240,
    UA_XOR_RF_IR210_A,
    UA__242,
    UA__243,
    UA_OR_RF_IR210_A,
    UA__245,
    UA__246,
    UA_AND_A_RF_IR210,
    UA__248,
    UA__249,
    UA_XOR_A_RF_IR210,
    UA__24B,
    UA__24C,
    UA_OR_A_RF_IR210,
    UA__24E,
    UA__24F,
    UA_CMPBNB_RF_IR210_A,
    UA__251,
    UA__252,
    UA_CMPB_RF_IR210_A,
    UA__254,
    UA__255,
    UA_CMPNZ_RF_IR210_A,
    UA__257,
    UA__258,
    UA_CMPZ_RF_IR210_A,
    UA__25A,
    UA__25B,
    UA_CMPBNB_A_RF_IR210,
    UA__25D,
    UA__25E,
    UA_CMPB_A_RF_IR210,
    UA__260,
    UA__261,
    UA_BITNZ_A_RF_IR210,
    UA__263,
    UA__264,
    UA_BITZ_A_RF_IR210,
    UA__266,
    UA__267,
    UA_CMPNZ_A_RF_IR210,
    UA__269,
    UA__26A,
    UA_CMPZ_A_RF_IR210,
    UA__26C,
    UA__26D,
    UA_ADDNC_RF_IR210_IMM,
    UA__26F,
    UA__270,
    UA__271,
    UA_SUBNB_RF_IR210_IMM,
    UA__273,
    UA__274,
    UA__275,
    UA_ADD_RF_IR210_IMM,
    UA__277,
    UA__278,
    UA__279,
    UA_ADC_RF_IR210_IMM,
    UA__27B,
    UA__27C,
    UA__27D,
    UA_SUB_RF_IR210_IMM,
    UA__27F,
    UA__280,
    UA__281,
    UA_SBB_RF_IR210_IMM,
    UA__283,
    UA__284,
    UA__285,
    UA_AND_RF_IR210_IMM,
    UA__287,
    UA__288,
    UA__289,
    UA_XOR_RF_IR210_IMM,
    UA__28B,
    UA__28C,
    UA__28D,
    UA_OR_RF_IR210_IMM,
    UA__28F,
    UA__290,
    UA__291,
    UA_ADDNC_SPR_IR2_IMM,
    UA__293,
    UA__294,
    UA__295,
    UA_SUBNB_SPR_IR2_IMM,
    UA__297,
    UA__298,
    UA__299,
    UA_ADD_SPR_IR2_IMM,
    UA__29B,
    UA__29C,
    UA__29D,
    UA_ADC_SPR_IR2_IMM,
    UA__29F,
    UA__2A0,
    UA__2A1,
    UA_SUB_SPR_IR2_IMM,
    UA__2A3,
    UA__2A4,
    UA__2A5,
    UA_SBB_SPR_IR2_IMM,
    UA__2A7,
    UA__2A8,
    UA__2A9,
    UA_AND_SPR_IR2_IMM,
    UA__2AB,
    UA__2AC,
    UA__2AD,
    UA_XOR_SPR_IR2_IMM,
    UA__2AF,
    UA__2B0,
    UA__2B1,
    UA_OR_SPR_IR2_IMM,
    UA__2B3,
    UA__2B4,
    UA__2B5,
    UA_CMPBNB_RF_IR210_IMM,
    UA__2B7,
    UA__2B8,
    UA__2B9,
    UA_CMPB_RF_IR210_IMM,
    UA__2BB,
    UA__2BC,
    UA__2BD,
    UA_BITNZ_RF_IR210_IMM,
    UA__2BF,
    UA__2C0,
    UA__2C1,
    UA_BITZ_RF_IR210_IMM,
    UA__2C3,
    UA__2C4,
    UA__2C5,
    UA_CMPNZ_RF_IR210_IMM,
    UA__2C7,
    UA__2C8,
    UA__2C9,
    UA_CMPZ_RF_IR210_IMM,
    UA__2CB,
    UA__2CC,
    UA__2CD,
    UA_CMPBNB_SPR_IR2_IMM,
    UA__2CF,
    UA__2D0,
    UA__2D1,
    UA_CMPB_SPR_IR2_IMM,
    UA__2D3,
    UA__2D4,
    UA__2D5,
    UA_BITNZ_SPR_IR2_IMM,
    UA__2D7,
    UA__2D8,
    UA__2D9,
    UA_BITZ_SPR_IR2_IMM,
    UA__2DB,
    UA__2DC,
    UA__2DD,
    UA_CMPNZ_SPR_IR2_IMM,
    UA__2DF,
    UA__2E0,
    UA__2E1,
    UA_CMPZ_SPR_IR2_IMM,
    UA__2E3,
    UA__2E4,
    UA__2E5,
    UA_LD_IR210_ABS,
    UA__2E7,
    UA__2E8,
    UA__2E9,
    UA__2EA,
    UA__2EB,
    UA__2EC,
    UA__2ED,
    UA__2EE,
    UA_LSPD,
    UA__2F0,
    UA__2F1,
    UA__2F2,
    UA__2F3,
    UA__2F4,
    UA__2F5,
    UA__2F6,
    UA__2F7,
    UA__2F8,
    UA__2F9,
    UA__2FA,
    UA_LBCD,
    UA__2FC,
    UA__2FD,
    UA__2FE,
    UA__2FF,
    UA__300,
    UA__301,
    UA__302,
    UA__303,
    UA__304,
    UA__305,
    UA__306,
    UA_LDED,
    UA__308,
    UA__309,
    UA__30A,
    UA__30B,
    UA__30C,
    UA__30D,
    UA__30E,
    UA__30F,
    UA__310,
    UA__311,
    UA__312,
    UA_LHLD,
    UA__314,
    UA__315,
    UA__316,
    UA__317,
    UA__318,
    UA__319,
    UA__31A,
    UA__31B,
    UA__31C,
    UA__31D,
    UA__31E,
    UA_ST_IR210_ABS,
    UA__320,
    UA__321,
    UA__322,
    UA__323,
    UA__324,
    UA__325,
    UA__326,
    UA__327,
    UA_SSPD,
    UA__329,
    UA__32A,
    UA__32B,
    UA__32C,
    UA__32D,
    UA__32E,
    UA__32F,
    UA__330,
    UA__331,
    UA__332,
    UA__333,
    UA_SBCD,
    UA__335,
    UA__336,
    UA__337,
    UA__338,
    UA__339,
    UA__33A,
    UA__33B,
    UA__33C,
    UA__33D,
    UA__33E,
    UA__33F,
    UA_SDED,
    UA__341,
    UA__342,
    UA__343,
    UA__344,
    UA__345,
    UA__346,
    UA__347,
    UA__348,
    UA__349,
    UA__34A,
    UA__34B,
    UA_SHLD,
    UA__34D,
    UA__34E,
    UA__34F,
    UA__350,
    UA__351,
    UA__352,
    UA__353,
    UA__354,
    UA__355,
    UA__356,
    UA__357,
    UA_ADDNC_A_IND,
    UA__359,
    UA__35A,
    UA__35B,
    UA_SUBNB_A_IND,
    UA__35D,
    UA__35E,
    UA__35F,
    UA_ADD_A_IND,
    UA__361,
    UA__362,
    UA__363,
    UA_ADC_A_IND,
    UA__365,
    UA__366,
    UA__367,
    UA_SUB_A_IND,
    UA__369,
    UA__36A,
    UA__36B,
    UA_SBB_A_IND,
    UA__36D,
    UA__36E,
    UA__36F,
    UA_AND_A_IND,
    UA__371,
    UA__372,
    UA__373,
    UA_XOR_A_IND,
    UA__375,
    UA__376,
    UA__377,
    UA_OR_A_IND,
    UA__379,
    UA__37A,
    UA__37B,
    UA_CMPBNB_A_IND,
    UA__37D,
    UA__37E,
    UA__37F,
    UA_CMPB_A_IND,
    UA__381,
    UA__382,
    UA__383,
    UA_BITNZ_A_IND,
    UA__385,
    UA__386,
    UA__387,
    UA_BITZ_A_IND,
    UA__389,
    UA__38A,
    UA__38B,
    UA_CMPNZ_A_IND,
    UA__38D,
    UA__38E,
    UA__38F,
    UA_CMPZ_A_IND,
    UA__391,
    UA__392,
    UA__393,
    UA_ADDNC_A_WA,
    UA__395,
    UA__396,
    UA__397,
    UA__398,
    UA__399,
    UA__39A,
    UA_SUBNB_A_WA,
    UA__39C,
    UA__39D,
    UA__39E,
    UA__39F,
    UA__3A0,
    UA__3A1,
    UA_ADD_A_WA,
    UA__3A3,
    UA__3A4,
    UA__3A5,
    UA__3A6,
    UA__3A7,
    UA__3A8,
    UA_ADC_A_WA,
    UA__3AA,
    UA__3AB,
    UA__3AC,
    UA__3AD,
    UA__3AE,
    UA__3AF,
    UA_SUB_A_WA,
    UA__3B1,
    UA__3B2,
    UA__3B3,
    UA__3B4,
    UA__3B5,
    UA__3B6,
    UA_SBB_A_WA,
    UA__3B8,
    UA__3B9,
    UA__3BA,
    UA__3BB,
    UA__3BC,
    UA__3BD,
    UA_AND_A_WA,
    UA__3BF,
    UA__3C0,
    UA__3C1,
    UA__3C2,
    UA__3C3,
    UA__3C4,
    UA_XOR_A_WA,
    UA__3C6,
    UA__3C7,
    UA__3C8,
    UA__3C9,
    UA__3CA,
    UA__3CB,
    UA_OR_A_WA,
    UA__3CD,
    UA__3CE,
    UA__3CF,
    UA__3D0,
    UA__3D1,
    UA__3D2,
    UA_CMPBNB_A_WA,
    UA__3D4,
    UA__3D5,
    UA__3D6,
    UA__3D7,
    UA__3D8,
    UA__3D9,
    UA_CMPB_A_WA,
    UA__3DB,
    UA__3DC,
    UA__3DD,
    UA__3DE,
    UA__3DF,
    UA__3E0,
    UA_BITNZ_A_WA,
    UA__3E2,
    UA__3E3,
    UA__3E4,
    UA__3E5,
    UA__3E6,
    UA__3E7,
    UA_BITZ_A_WA,
    UA__3E9,
    UA__3EA,
    UA__3EB,
    UA__3EC,
    UA__3ED,
    UA__3EE,
    UA_CMPNZ_A_WA,
    UA__3F0,
    UA__3F1,
    UA__3F2,
    UA__3F3,
    UA__3F4,
    UA__3F5,
    UA_CMPZ_A_WA,
    UA__3F7,
    UA__3F8,
    UA__3F9,
    UA__3FA,
    UA__3FB,
    UA__3FC
} e_uaddr;    // ucode address

typedef reg [7:0] t_naddr;    // ncode address

typedef enum reg [1:0]
{
    UBM_ADV,
    UBM_END,
    UBM_DA
} e_ubm;    // branch mode

typedef enum reg [1:0]
{
    UTX_T1,
    UTX_T2,
    UTX_T3,
    UTX_T4
} e_mcy;    // machine cycle

typedef enum reg [3:0]
{
    URFS_V,
    URFS_A,
    URFS_B,
    URFS_C,
    URFS_D,
    URFS_E,
    URFS_H,
    URFS_L,
    URFS_PSW,
    URFS_SPL,
    URFS_SPH,
    URFS_PCL,
    URFS_PCH,
    URFS_IR210,
    URFS_W
} e_urfs;    // register file select

typedef enum reg [2:0]
{
    UIDBS_0,
    UIDBS_RF,
    UIDBS_DB,
    UIDBS_CO,
    UIDBS_SPR,
    UIDBS_SDG
} e_idbs;    // idb select

typedef enum reg [3:0]
{
    ULTS_NONE,
    ULTS_RF,
    ULTS_DOR,
    ULTS_AI,
    ULTS_BI,
    ULTS_IE,
    ULTS_SPR,
    ULTS_PSW_CY
} e_lts;    // load target select

typedef enum reg [3:0]
{
    UABS_PC,
    UABS_SP,
    UABS_BC,
    UABS_DE,
    UABS_HL,
    UABS_VW,
    UABS_IDB_W,
    UABS_IR210,
    UABS_AOR,
    UABS_NABI
} e_abs;    // ab select

typedef enum reg [3:0]
{
    USPR_PA,
    USPR_PB,
    USPR_PC,
    USPR_MK,
    USPR_MB,
    USPR_MC,
    USPR_TM0,
    USPR_TM1,
    USPR_S,
    USPR_TMM
} e_spr;    // special register

typedef enum reg [0:0]
{
    USRS_IR2,
    USRS_IR3
} e_sprs;    // special register select

typedef enum reg [2:0]
{
    USDGS_JRL,
    USDGS_JRH,
    USDGS_CALF,
    USDGS_CALT,
    USDGS_INTVA,
    USDGS_BIT
} e_sdgs;    // special data generator select

typedef enum reg [3:0]
{
    UAO_NOP,
    UAO_SUM,
    UAO_SUB,
    UAO_INC,
    UAO_DEC,
    UAO_OR,
    UAO_AND,
    UAO_EOR,
    UAO_LSL,
    UAO_ROL,
    UAO_LSR,
    UAO_ROR,
    UAO_DIL,
    UAO_DIH,
    UAO_DIS
} e_aluop;    // ALU operation

typedef enum reg [1:0]
{
    UCIS_0,
    UCIS_1,
    UCIS_CCO,
    UCIS_PSW_CY
} e_cis;    // ALU carry in select

typedef enum reg [3:0]
{
    USKS_PSW_SK,
    USKS_1,
    USKS_C,
    USKS_NC,
    USKS_Z,
    USKS_NZ,
    USKS_I,
    USKS_NI,
    USKS_0,
    USKS_PSW_C,
    USKS_PSW_NC,
    USKS_PSW_Z,
    USKS_PSW_NZ
} e_sks;    // SKip flag source

typedef struct packed
{
    e_uaddr uaddr;    // microcode entry point
    reg [0:0] m1_overlap;    // New M1 starts immediately
    reg [1:0] skipn;    // Number of operands to skip when ins. is skipped
} s_ird;

typedef struct packed
{
    t_naddr naddr;    // nanocode address
    e_ubm bm;    // branch mode
    reg [0:0] m1;    // Fetch next opcode (start M1)
} s_uc;

typedef struct packed
{
    reg [2:0] idx;    // general-purpose data
    e_urfs rfos;    // register file output select -> idb
    e_urfs rfts;    // register file target select
    e_idbs idbs;    // idb select
    e_lts lts;    // load target select
    e_abs abs;    // ab select
    e_abs abits;    // abi target select
    reg [0:0] pc_inc;    // increment PC
    reg [0:0] ab_inc;    // increment ab
    reg [0:0] ab_dec;    // decrement ab
    reg [0:0] aout;    // ab -> AOR
    reg [0:0] load;    // assert RDB (read operation)
    reg [0:0] store;    // dor -> DB
    e_aluop aluop;    // ALU operation
    e_cis cis;    // ALU carry in select
    reg [0:0] bi0;    // Zero BI
    reg [0:0] bin;    // Negate BI
    reg [0:0] pswz;    // (CO == 0) -> PSW.Z
    reg [0:0] pswcy;    // CCO -> PSW.CY
    reg [0:0] pswhc;    // CHO -> PSW.HC
    e_sks pswsk;    // PSW.SK source
    e_sprs sprs;    // special register select
    e_sdgs sdgs;    // special data generator select
    reg [0:0] daa;    // decimal adjust const -> BI
    reg [0:0] rpir;    // IR[2:0] selects reg. pair and inc/dec
} s_nc;

