s_nc nrom [194];
initial begin
  nrom[   0] = 53'b00000000000000000000000000000000000000000000000000000;
  nrom[   1] = 53'b00000000000000000000000000100100000000000000000000000;
  nrom[   2] = 53'b00000000000000000000000000000010000000000000000000000;
  nrom[   3] = 53'b00000000000000000000000000000001000000000000000000000;
  nrom[   4] = 53'b00011010001001000100000000000000000000000000000000000;
  nrom[   5] = 53'b00000011101001000100000000000000000000000000000000000;
  nrom[   6] = 53'b00000001101010000100000000000000000000000000000000000;
  nrom[   7] = 53'b00000001110010000100000000000000000000000000000000000;
  nrom[   8] = 53'b00000000000000000001010000000100000000000000000000000;
  nrom[   9] = 53'b00000000001010000100000000000000000000000000000000000;
  nrom[  10] = 53'b00000001001010000100000000000000000000000000000000000;
  nrom[  11] = 53'b00000001010010000100000000000000000000000000000000000;
  nrom[  12] = 53'b00000000011010000100000000000000000000000000000000000;
  nrom[  13] = 53'b00000000010010000100000000000000000000000000000000000;
  nrom[  14] = 53'b00000000101010000100000000000000000000000000000000000;
  nrom[  15] = 53'b00000000100010000100000000000000000000000000000000000;
  nrom[  16] = 53'b00000000111010000100000000000000000000000000000000000;
  nrom[  17] = 53'b00000000110010000100000000000000000000000000000000000;
  nrom[  18] = 53'b00000000000000000001110111000100000000000000000000001;
  nrom[  19] = 53'b00000010000001001001110111000100000000000000000000001;
  nrom[  20] = 53'b00011100000001001001110111000100000000000000000000001;
  nrom[  21] = 53'b00000010000001001001010000000100000000000000000000000;
  nrom[  22] = 53'b00000000000010001100000000000000000100100000000000000;
  nrom[  23] = 53'b00000000000011001001010000000100000000000000000000000;
  nrom[  24] = 53'b00010110000001001100000000000000000000000000000000000;
  nrom[  25] = 53'b00000010000001010000000000000000000101000000000000000;
  nrom[  26] = 53'b00000001110011000100000000000000000000000000000000000;
  nrom[  27] = 53'b00011000000001001100000000000000000110100000000000000;
  nrom[  28] = 53'b00000000000011000001100000000100000000000000000000000;
  nrom[  29] = 53'b00000000011010000110000000000000000000000000000000000;
  nrom[  30] = 53'b00000000000000000010010000010100000000000000000000000;
  nrom[  31] = 53'b00000000000000000001000000000100000000000000000000000;
  nrom[  32] = 53'b00000000000000000001000100010010000000000000000000000;
  nrom[  33] = 53'b00011100000001001000110000000100000000000000000000000;
  nrom[  34] = 53'b00000000000000000000110011010001000000000000000000000;
  nrom[  35] = 53'b00000110000001001100000000000000010000000000000000000;
  nrom[  36] = 53'b00000000011011000100000000000000000000000000000000000;
  nrom[  37] = 53'b00000000000000000000000000001000000000000000010000000;
  nrom[  38] = 53'b00000000000010001100000000000000000000000000000000000;
  nrom[  39] = 53'b00000000000010010000000000000000011000000000000000000;
  nrom[  40] = 53'b00000000000000000000000000000000000000001000000000000;
  nrom[  41] = 53'b00000000000010010000000000000000010100000000000000000;
  nrom[  42] = 53'b00000010000001001100000000100100000000000000000000000;
  nrom[  43] = 53'b00000000001011000100000000000000000000001000000000000;
  nrom[  44] = 53'b00000000000010010000000000000000011100000000000000000;
  nrom[  45] = 53'b00000000000010010000000000000000001001010000000000000;
  nrom[  46] = 53'b00000000000000000000000000000000000000001110011000000;
  nrom[  47] = 53'b00000000000010010000000000000000001000010000000000000;
  nrom[  48] = 53'b00000000000000000000000000000000000000001110010000000;
  nrom[  49] = 53'b00000000000000000000000000000000000000001000101000000;
  nrom[  50] = 53'b00000000000000000000000000000000000000001000100000000;
  nrom[  51] = 53'b00000000000000000000000000000000000000001110101000000;
  nrom[  52] = 53'b00000000000000000000000000000000000000001110100000000;
  nrom[  53] = 53'b00000000000010010000000000000000000100000000000000000;
  nrom[  54] = 53'b00000000001011000100000000000000000000001110011000000;
  nrom[  55] = 53'b00000000000010010000000000000000001000010000000000000;
  nrom[  56] = 53'b00000000001011000100000000000000000000001110000000000;
  nrom[  57] = 53'b00000000000010010000000000000000000111000000000000000;
  nrom[  58] = 53'b00000000000010010000000000000000001011010000000000000;
  nrom[  59] = 53'b00000000000010001100000000000000001100000000000000000;
  nrom[  60] = 53'b00000000000000000000000000000000000000001010010000000;
  nrom[  61] = 53'b00000000000010001100000000000000010000000000000000000;
  nrom[  62] = 53'b00011010000001001100000000000000001100000000000000000;
  nrom[  63] = 53'b00000001101011000100000000000000000000001010010000000;
  nrom[  64] = 53'b00011010000001001100000000000000010000000000000000000;
  nrom[  65] = 53'b00000000000000000000010001010000000000000000000000000;
  nrom[  66] = 53'b00000000000000000000100010010000000000000000000000000;
  nrom[  67] = 53'b00000000000000000000110011010000000000000000000000000;
  nrom[  68] = 53'b00000000000000000001000100010000000000000000000000000;
  nrom[  69] = 53'b00000000000000000000010001001000000000000000000000000;
  nrom[  70] = 53'b00000000000000000000100010001000000000000000000000000;
  nrom[  71] = 53'b00000000000000000000110011001000000000000000000000000;
  nrom[  72] = 53'b00000000000000000001000100001000000000000000000000000;
  nrom[  73] = 53'b00000010000001001100000000000000000100000000000000010;
  nrom[  74] = 53'b00000000000101010000000000000000000000000000000000000;
  nrom[  75] = 53'b00000000000000000000000000000000000100000000000000000;
  nrom[  76] = 53'b00000001011011000100000000000000000000000000000000000;
  nrom[  77] = 53'b00011000000001001100000000000000000000000000000000000;
  nrom[  78] = 53'b00000000000101010000000000000000000000000000000000100;
  nrom[  79] = 53'b00000000000000000000000000000000000110000000000000000;
  nrom[  80] = 53'b00000001100011000100000000000000000000000000000000000;
  nrom[  81] = 53'b00010110000001001100000000000010000000000000000000000;
  nrom[  82] = 53'b00000000000010010000000000000000000100000000000000000;
  nrom[  83] = 53'b00011000000001001100000000000000000110100000000000000;
  nrom[  84] = 53'b00011000000001001100000000000000000110110000000000000;
  nrom[  85] = 53'b00000000000000000000000000000100000000000000000000000;
  nrom[  86] = 53'b00011101011001000100000000000010000000000000000000000;
  nrom[  87] = 53'b00000001100010000100000000000000000000000000000000000;
  nrom[  88] = 53'b00000000000000000000100000011100000000000000000000000;
  nrom[  89] = 53'b00000000000010001100010001001000000100100000000000000;
  nrom[  90] = 53'b00011000000001001000010000000100000000000000000000000;
  nrom[  91] = 53'b00010110000001001000010000000100000000000000000000000;
  nrom[  92] = 53'b00011101011001000100000000000001000000000000000000000;
  nrom[  93] = 53'b00000101100001000100000000000001000000000000000000000;
  nrom[  94] = 53'b00000111011001000100000000000001000000000000000000000;
  nrom[  95] = 53'b00000000000000000000000000100000000000000000000000000;
  nrom[  96] = 53'b00000001110010000100010001001000000000000000000000000;
  nrom[  97] = 53'b00000000000000000000000000001000000000000000000000000;
  nrom[  98] = 53'b00000001100101000100000000000010000000000000000001000;
  nrom[  99] = 53'b00000001011010000100000000000000000000000000000000000;
  nrom[ 100] = 53'b00000001110101000100000000000000000000000000000001100;
  nrom[ 101] = 53'b00000000000000000001100000000100000000000000000000000;
  nrom[ 102] = 53'b00100001110101000100000000000010000000000000000001100;
  nrom[ 103] = 53'b00010000000001001000010000000100000000000000000000000;
  nrom[ 104] = 53'b00000001100000000100000000000000000000000000000000000;
  nrom[ 105] = 53'b00000001011101000100000000000000000000000000000010000;
  nrom[ 106] = 53'b00000000000000000000000000000000000000000001000000000;
  nrom[ 107] = 53'b00000000000000000000010000000100000000000000000000000;
  nrom[ 108] = 53'b00000000000000000000010001010010000000000000000000000;
  nrom[ 109] = 53'b00000001100010000100000000000000000000000000001000000;
  nrom[ 110] = 53'b00000001000010000100000000000000000000000000000000000;
  nrom[ 111] = 53'b00000000000101010000000000000010000000000000000010100;
  nrom[ 112] = 53'b00000000000010001100000000000000011000000000000000000;
  nrom[ 113] = 53'b00000000000000000000000000000000000000000000101000000;
  nrom[ 114] = 53'b00000010000001001100000000000000000000000000000000000;
  nrom[ 115] = 53'b00000000000000000000000000000000100111000000000000000;
  nrom[ 116] = 53'b00000000001011000100000000000000000000000100000000000;
  nrom[ 117] = 53'b00000000000000000000000000000000101111000000000000000;
  nrom[ 118] = 53'b00000110000001001100000000000000000000000000000000000;
  nrom[ 119] = 53'b00000000011011000100000000000000000000000100000000000;
  nrom[ 120] = 53'b00000000000000000000000000000000100000000000000000000;
  nrom[ 121] = 53'b00000000000000000000000000000000101000000000000000000;
  nrom[ 122] = 53'b00000000000001001000010000000100000000000000000000000;
  nrom[ 123] = 53'b00000010000001001000010000000100000000000000000000000;
  nrom[ 124] = 53'b00000000000000000000010001010100000000000000000000000;
  nrom[ 125] = 53'b00000000000010000100000000000000000000000000000000000;
  nrom[ 126] = 53'b00000100000001001000010000000100000000000000000000000;
  nrom[ 127] = 53'b00000110000001001000010000000100000000000000000000000;
  nrom[ 128] = 53'b00001000000001001000010000000100000000000000000000000;
  nrom[ 129] = 53'b00001010000001001000010000000100000000000000000000000;
  nrom[ 130] = 53'b00001100000001001000010000000100000000000000000000000;
  nrom[ 131] = 53'b00001110000001001000010000000100000000000000000000000;
  nrom[ 132] = 53'b00000000000000000000000000000000000000000000110000000;
  nrom[ 133] = 53'b00000000000000000000000000000000000000000001001000000;
  nrom[ 134] = 53'b00000000000000000000000000000000000000000001011000000;
  nrom[ 135] = 53'b00000000000000000000000000000000000000000000111000000;
  nrom[ 136] = 53'b00000000000000000000000000000000000000000001010000000;
  nrom[ 137] = 53'b00000000000000000000000000000000000000000001100000000;
  nrom[ 138] = 53'b00100000000000010100000000000000000000000000000000000;
  nrom[ 139] = 53'b00000000000000010100000000000000000000000000000000000;
  nrom[ 140] = 53'b00000000000000011100000000000000000000000000000000000;
  nrom[ 141] = 53'b00100000000000011100000000000000000000000000000000000;
  nrom[ 142] = 53'b00011100000001001100000000000000111000000000000000000;
  nrom[ 143] = 53'b00000010000001001100000000000000110000000000000000000;
  nrom[ 144] = 53'b00011100000011001001000000000100000000000000000000000;
  nrom[ 145] = 53'b00011100000001001100000000000001110000000000000000000;
  nrom[ 146] = 53'b00000010000001001100000000000000110100000000000000000;
  nrom[ 147] = 53'b00000000001011000100000000000000000000000000000000000;
  nrom[ 148] = 53'b00011100000001001100000000000000110100000000000000000;
  nrom[ 149] = 53'b00000000000011001100000000000000111000000000000000000;
  nrom[ 150] = 53'b00000000001100000100000000000000000000000000000100000;
  nrom[ 151] = 53'b00000010000001011000000000000000000000000000000100000;
  nrom[ 152] = 53'b00011010000001001100000000000000000000000000000000000;
  nrom[ 153] = 53'b00000010000001010000000000000000000100000000000000000;
  nrom[ 154] = 53'b00000001101011000100000000000000000000001110011000000;
  nrom[ 155] = 53'b00000010000001010000000000000000001000010000000000000;
  nrom[ 156] = 53'b00000001101011000100000000000000000000001110000000000;
  nrom[ 157] = 53'b00000010000001010000000000000000000111000000000000000;
  nrom[ 158] = 53'b00000010000001010000000000000000001011010000000000000;
  nrom[ 159] = 53'b00011010000001010000000000000000000100000000000000000;
  nrom[ 160] = 53'b00011010000001010000000000000000001000010000000000000;
  nrom[ 161] = 53'b00011010000001010000000000000000000111000000000000000;
  nrom[ 162] = 53'b00011010000001010000000000000000001011010000000000000;
  nrom[ 163] = 53'b00000010000001010000000000000000011000000000000000000;
  nrom[ 164] = 53'b00000001101011000100000000000000000000001000000000000;
  nrom[ 165] = 53'b00000010000001010000000000000000011100000000000000000;
  nrom[ 166] = 53'b00000010000001010000000000000000010100000000000000000;
  nrom[ 167] = 53'b00011010000001010000000000000000011000000000000000000;
  nrom[ 168] = 53'b00011010000001010000000000000000011100000000000000000;
  nrom[ 169] = 53'b00011010000001010000000000000000010100000000000000000;
  nrom[ 170] = 53'b00000010000001010000000000000000001001010000000000000;
  nrom[ 171] = 53'b00000010000001010000000000000000001000010000000000000;
  nrom[ 172] = 53'b00011010000001010000000000000000001001010000000000000;
  nrom[ 173] = 53'b00011010000001010000000000000000001000010000000000000;
  nrom[ 174] = 53'b00011010000001001100000000100100000000000000000000000;
  nrom[ 175] = 53'b00000000000100001100000000100100000000000000000000000;
  nrom[ 176] = 53'b00000000000011011000000000000000000000001110011000000;
  nrom[ 177] = 53'b00000000000011011000000000000000000000001110000000000;
  nrom[ 178] = 53'b00000000000011011000000000000000000000001000000000000;
  nrom[ 179] = 53'b00000001001010000110000000000000000000000000000000000;
  nrom[ 180] = 53'b00000000101010000110000000000000000000000000000000000;
  nrom[ 181] = 53'b00000000111010000110000000000000000000000000000000000;
  nrom[ 182] = 53'b00011010000001001000000000000010000000000000000000000;
  nrom[ 183] = 53'b00010010000001001000000000000010000000000000000000000;
  nrom[ 184] = 53'b00000000000000000010000000000000000000000000000000000;
  nrom[ 185] = 53'b00010100000001001010010000010100000000000000000000000;
  nrom[ 186] = 53'b00000110000001001000000000000010000000000000000000000;
  nrom[ 187] = 53'b00000100000001001010010000010100000000000000000000000;
  nrom[ 188] = 53'b00001010000001001000000000000010000000000000000000000;
  nrom[ 189] = 53'b00001000000001001010010000010100000000000000000000000;
  nrom[ 190] = 53'b00001110000001001000000000000010000000000000000000000;
  nrom[ 191] = 53'b00001100000001001010010000010100000000000000000000000;
  nrom[ 192] = 53'b00000010000001001100000000000010000000000000000000000;
  nrom[ 193] = 53'b00000010000001001101010000000100000000000000000000000;
end
